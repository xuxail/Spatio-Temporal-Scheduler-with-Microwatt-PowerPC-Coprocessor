VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openframe_project_wrapper
  CLASS BLOCK ;
  FOREIGN openframe_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3166.630 BY 4766.630 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 306.190 3168.630 306.830 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3222.190 3168.630 3222.830 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3447.190 3168.630 3447.830 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3672.190 3168.630 3672.830 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4118.190 3168.630 4118.830 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4564.190 3168.630 4564.830 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2981.800 4766.350 2982.440 4768.630 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.800 4766.350 2473.440 4768.630 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.800 4766.350 2216.440 4768.630 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.800 4766.350 1771.440 4768.630 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.800 4766.350 1262.440 4768.630 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 532.190 3168.630 532.830 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.800 4766.350 1004.440 4768.630 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.800 4766.350 747.440 4768.630 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.800 4766.350 490.440 4768.630 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.800 4766.350 233.440 4768.630 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4622.800 0.300 4623.440 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3773.800 0.300 3774.440 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3557.800 0.300 3558.440 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3341.800 0.300 3342.440 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3125.800 0.300 3126.440 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2909.800 0.300 2910.440 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 757.190 3168.630 757.830 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2693.800 0.300 2694.440 ;
    END
  END analog_io[30]
  PIN analog_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2477.800 0.300 2478.440 ;
    END
  END analog_io[31]
  PIN analog_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1839.800 0.300 1840.440 ;
    END
  END analog_io[32]
  PIN analog_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1623.800 0.300 1624.440 ;
    END
  END analog_io[33]
  PIN analog_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1407.800 0.300 1408.440 ;
    END
  END analog_io[34]
  PIN analog_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1191.800 0.300 1192.440 ;
    END
  END analog_io[35]
  PIN analog_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 975.800 0.300 976.440 ;
    END
  END analog_io[36]
  PIN analog_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 759.800 0.300 760.440 ;
    END
  END analog_io[37]
  PIN analog_io[38]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.190 -2.000 738.830 0.280 ;
    END
  END analog_io[38]
  PIN analog_io[39]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.190 -2.000 1281.830 0.280 ;
    END
  END analog_io[39]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 983.190 3168.630 983.830 ;
    END
  END analog_io[3]
  PIN analog_io[40]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.190 -2.000 1555.830 0.280 ;
    END
  END analog_io[40]
  PIN analog_io[41]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.190 -2.000 1829.830 0.280 ;
    END
  END analog_io[41]
  PIN analog_io[42]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.190 -2.000 2103.830 0.280 ;
    END
  END analog_io[42]
  PIN analog_io[43]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.190 -2.000 2377.830 0.280 ;
    END
  END analog_io[43]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1208.190 3168.630 1208.830 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1433.190 3168.630 1433.830 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1659.190 3168.630 1659.830 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2545.190 3168.630 2545.830 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2771.190 3168.630 2771.830 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2996.190 3168.630 2996.830 ;
    END
  END analog_io[9]
  PIN analog_noesd_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 315.175 3168.630 316.245 ;
    END
  END analog_noesd_io[0]
  PIN analog_noesd_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3231.175 3168.630 3232.245 ;
    END
  END analog_noesd_io[10]
  PIN analog_noesd_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3456.175 3168.630 3457.245 ;
    END
  END analog_noesd_io[11]
  PIN analog_noesd_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3681.175 3168.630 3682.245 ;
    END
  END analog_noesd_io[12]
  PIN analog_noesd_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4127.175 3168.630 4128.245 ;
    END
  END analog_noesd_io[13]
  PIN analog_noesd_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4573.175 3168.630 4574.245 ;
    END
  END analog_noesd_io[14]
  PIN analog_noesd_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2972.385 4766.350 2973.455 4768.630 ;
    END
  END analog_noesd_io[15]
  PIN analog_noesd_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.385 4766.350 2464.455 4768.630 ;
    END
  END analog_noesd_io[16]
  PIN analog_noesd_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.385 4766.350 2207.455 4768.630 ;
    END
  END analog_noesd_io[17]
  PIN analog_noesd_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.385 4766.350 1762.455 4768.630 ;
    END
  END analog_noesd_io[18]
  PIN analog_noesd_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.385 4766.350 1253.455 4768.630 ;
    END
  END analog_noesd_io[19]
  PIN analog_noesd_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 541.175 3168.630 542.245 ;
    END
  END analog_noesd_io[1]
  PIN analog_noesd_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.385 4766.350 995.455 4768.630 ;
    END
  END analog_noesd_io[20]
  PIN analog_noesd_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.385 4766.350 738.455 4768.630 ;
    END
  END analog_noesd_io[21]
  PIN analog_noesd_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.385 4766.350 481.455 4768.630 ;
    END
  END analog_noesd_io[22]
  PIN analog_noesd_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.385 4766.350 224.455 4768.630 ;
    END
  END analog_noesd_io[23]
  PIN analog_noesd_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4613.385 0.300 4614.455 ;
    END
  END analog_noesd_io[24]
  PIN analog_noesd_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3764.385 0.300 3765.455 ;
    END
  END analog_noesd_io[25]
  PIN analog_noesd_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3548.385 0.300 3549.455 ;
    END
  END analog_noesd_io[26]
  PIN analog_noesd_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3332.385 0.300 3333.455 ;
    END
  END analog_noesd_io[27]
  PIN analog_noesd_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3116.385 0.300 3117.455 ;
    END
  END analog_noesd_io[28]
  PIN analog_noesd_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2900.385 0.300 2901.455 ;
    END
  END analog_noesd_io[29]
  PIN analog_noesd_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 766.175 3168.630 767.245 ;
    END
  END analog_noesd_io[2]
  PIN analog_noesd_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2684.385 0.300 2685.455 ;
    END
  END analog_noesd_io[30]
  PIN analog_noesd_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2468.385 0.300 2469.455 ;
    END
  END analog_noesd_io[31]
  PIN analog_noesd_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1830.385 0.300 1831.455 ;
    END
  END analog_noesd_io[32]
  PIN analog_noesd_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1614.385 0.300 1615.455 ;
    END
  END analog_noesd_io[33]
  PIN analog_noesd_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1398.385 0.300 1399.455 ;
    END
  END analog_noesd_io[34]
  PIN analog_noesd_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1182.385 0.300 1183.455 ;
    END
  END analog_noesd_io[35]
  PIN analog_noesd_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 966.385 0.300 967.455 ;
    END
  END analog_noesd_io[36]
  PIN analog_noesd_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 750.385 0.300 751.455 ;
    END
  END analog_noesd_io[37]
  PIN analog_noesd_io[38]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.175 -2.000 748.245 0.280 ;
    END
  END analog_noesd_io[38]
  PIN analog_noesd_io[39]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.175 -2.000 1291.245 0.280 ;
    END
  END analog_noesd_io[39]
  PIN analog_noesd_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 992.175 3168.630 993.245 ;
    END
  END analog_noesd_io[3]
  PIN analog_noesd_io[40]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.175 -2.000 1565.245 0.280 ;
    END
  END analog_noesd_io[40]
  PIN analog_noesd_io[41]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.175 -2.000 1839.245 0.280 ;
    END
  END analog_noesd_io[41]
  PIN analog_noesd_io[42]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.175 -2.000 2113.245 0.280 ;
    END
  END analog_noesd_io[42]
  PIN analog_noesd_io[43]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.175 -2.000 2387.245 0.280 ;
    END
  END analog_noesd_io[43]
  PIN analog_noesd_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1217.175 3168.630 1218.245 ;
    END
  END analog_noesd_io[4]
  PIN analog_noesd_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1442.175 3168.630 1443.245 ;
    END
  END analog_noesd_io[5]
  PIN analog_noesd_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1668.175 3168.630 1669.245 ;
    END
  END analog_noesd_io[6]
  PIN analog_noesd_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2554.175 3168.630 2555.245 ;
    END
  END analog_noesd_io[7]
  PIN analog_noesd_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2780.175 3168.630 2781.245 ;
    END
  END analog_noesd_io[8]
  PIN analog_noesd_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3005.175 3168.630 3006.245 ;
    END
  END analog_noesd_io[9]
  PIN gpio_analog_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 318.300 3168.630 318.650 ;
    END
  END gpio_analog_en[0]
  PIN gpio_analog_en[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3234.300 3168.630 3234.650 ;
    END
  END gpio_analog_en[10]
  PIN gpio_analog_en[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3459.300 3168.630 3459.650 ;
    END
  END gpio_analog_en[11]
  PIN gpio_analog_en[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3684.300 3168.630 3684.650 ;
    END
  END gpio_analog_en[12]
  PIN gpio_analog_en[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4130.300 3168.630 4130.650 ;
    END
  END gpio_analog_en[13]
  PIN gpio_analog_en[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4576.300 3168.630 4576.650 ;
    END
  END gpio_analog_en[14]
  PIN gpio_analog_en[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2970.020 4766.350 2970.300 4768.630 ;
    END
  END gpio_analog_en[15]
  PIN gpio_analog_en[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.020 4766.350 2461.300 4768.630 ;
    END
  END gpio_analog_en[16]
  PIN gpio_analog_en[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.020 4766.350 2204.300 4768.630 ;
    END
  END gpio_analog_en[17]
  PIN gpio_analog_en[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.020 4766.350 1759.300 4768.630 ;
    END
  END gpio_analog_en[18]
  PIN gpio_analog_en[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.020 4766.350 1250.300 4768.630 ;
    END
  END gpio_analog_en[19]
  PIN gpio_analog_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 544.300 3168.630 544.650 ;
    END
  END gpio_analog_en[1]
  PIN gpio_analog_en[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.020 4766.350 992.300 4768.630 ;
    END
  END gpio_analog_en[20]
  PIN gpio_analog_en[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.020 4766.350 735.300 4768.630 ;
    END
  END gpio_analog_en[21]
  PIN gpio_analog_en[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.020 4766.350 478.300 4768.630 ;
    END
  END gpio_analog_en[22]
  PIN gpio_analog_en[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.020 4766.350 221.300 4768.630 ;
    END
  END gpio_analog_en[23]
  PIN gpio_analog_en[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4610.980 0.300 4611.330 ;
    END
  END gpio_analog_en[24]
  PIN gpio_analog_en[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3761.980 0.300 3762.330 ;
    END
  END gpio_analog_en[25]
  PIN gpio_analog_en[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3545.980 0.300 3546.330 ;
    END
  END gpio_analog_en[26]
  PIN gpio_analog_en[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3329.980 0.300 3330.330 ;
    END
  END gpio_analog_en[27]
  PIN gpio_analog_en[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3113.980 0.300 3114.330 ;
    END
  END gpio_analog_en[28]
  PIN gpio_analog_en[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2897.980 0.300 2898.330 ;
    END
  END gpio_analog_en[29]
  PIN gpio_analog_en[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 769.300 3168.630 769.650 ;
    END
  END gpio_analog_en[2]
  PIN gpio_analog_en[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2681.980 0.300 2682.330 ;
    END
  END gpio_analog_en[30]
  PIN gpio_analog_en[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2465.980 0.300 2466.330 ;
    END
  END gpio_analog_en[31]
  PIN gpio_analog_en[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1827.980 0.300 1828.330 ;
    END
  END gpio_analog_en[32]
  PIN gpio_analog_en[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1611.980 0.300 1612.330 ;
    END
  END gpio_analog_en[33]
  PIN gpio_analog_en[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1395.980 0.300 1396.330 ;
    END
  END gpio_analog_en[34]
  PIN gpio_analog_en[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1179.980 0.300 1180.330 ;
    END
  END gpio_analog_en[35]
  PIN gpio_analog_en[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 963.980 0.300 964.330 ;
    END
  END gpio_analog_en[36]
  PIN gpio_analog_en[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 747.980 0.300 748.330 ;
    END
  END gpio_analog_en[37]
  PIN gpio_analog_en[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.330 -2.000 750.610 0.280 ;
    END
  END gpio_analog_en[38]
  PIN gpio_analog_en[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.330 -2.000 1293.610 0.280 ;
    END
  END gpio_analog_en[39]
  PIN gpio_analog_en[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 995.300 3168.630 995.650 ;
    END
  END gpio_analog_en[3]
  PIN gpio_analog_en[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.330 -2.000 1567.610 0.280 ;
    END
  END gpio_analog_en[40]
  PIN gpio_analog_en[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.330 -2.000 1841.610 0.280 ;
    END
  END gpio_analog_en[41]
  PIN gpio_analog_en[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.330 -2.000 2115.610 0.280 ;
    END
  END gpio_analog_en[42]
  PIN gpio_analog_en[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.330 -2.000 2389.610 0.280 ;
    END
  END gpio_analog_en[43]
  PIN gpio_analog_en[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1220.300 3168.630 1220.650 ;
    END
  END gpio_analog_en[4]
  PIN gpio_analog_en[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1445.300 3168.630 1445.650 ;
    END
  END gpio_analog_en[5]
  PIN gpio_analog_en[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1671.300 3168.630 1671.650 ;
    END
  END gpio_analog_en[6]
  PIN gpio_analog_en[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2557.300 3168.630 2557.650 ;
    END
  END gpio_analog_en[7]
  PIN gpio_analog_en[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2783.300 3168.630 2783.650 ;
    END
  END gpio_analog_en[8]
  PIN gpio_analog_en[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3008.300 3168.630 3008.650 ;
    END
  END gpio_analog_en[9]
  PIN gpio_analog_pol[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 324.740 3168.630 325.090 ;
    END
  END gpio_analog_pol[0]
  PIN gpio_analog_pol[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3240.740 3168.630 3241.090 ;
    END
  END gpio_analog_pol[10]
  PIN gpio_analog_pol[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3465.740 3168.630 3466.090 ;
    END
  END gpio_analog_pol[11]
  PIN gpio_analog_pol[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3690.740 3168.630 3691.090 ;
    END
  END gpio_analog_pol[12]
  PIN gpio_analog_pol[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4136.740 3168.630 4137.090 ;
    END
  END gpio_analog_pol[13]
  PIN gpio_analog_pol[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4582.740 3168.630 4583.090 ;
    END
  END gpio_analog_pol[14]
  PIN gpio_analog_pol[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2963.580 4766.350 2963.860 4768.630 ;
    END
  END gpio_analog_pol[15]
  PIN gpio_analog_pol[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.580 4766.350 2454.860 4768.630 ;
    END
  END gpio_analog_pol[16]
  PIN gpio_analog_pol[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.580 4766.350 2197.860 4768.630 ;
    END
  END gpio_analog_pol[17]
  PIN gpio_analog_pol[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.580 4766.350 1752.860 4768.630 ;
    END
  END gpio_analog_pol[18]
  PIN gpio_analog_pol[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.580 4766.350 1243.860 4768.630 ;
    END
  END gpio_analog_pol[19]
  PIN gpio_analog_pol[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 550.740 3168.630 551.090 ;
    END
  END gpio_analog_pol[1]
  PIN gpio_analog_pol[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.580 4766.350 985.860 4768.630 ;
    END
  END gpio_analog_pol[20]
  PIN gpio_analog_pol[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.580 4766.350 728.860 4768.630 ;
    END
  END gpio_analog_pol[21]
  PIN gpio_analog_pol[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.580 4766.350 471.860 4768.630 ;
    END
  END gpio_analog_pol[22]
  PIN gpio_analog_pol[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.580 4766.350 214.860 4768.630 ;
    END
  END gpio_analog_pol[23]
  PIN gpio_analog_pol[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4604.540 0.300 4604.890 ;
    END
  END gpio_analog_pol[24]
  PIN gpio_analog_pol[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3755.540 0.300 3755.890 ;
    END
  END gpio_analog_pol[25]
  PIN gpio_analog_pol[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3539.540 0.300 3539.890 ;
    END
  END gpio_analog_pol[26]
  PIN gpio_analog_pol[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3323.540 0.300 3323.890 ;
    END
  END gpio_analog_pol[27]
  PIN gpio_analog_pol[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3107.540 0.300 3107.890 ;
    END
  END gpio_analog_pol[28]
  PIN gpio_analog_pol[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2891.540 0.300 2891.890 ;
    END
  END gpio_analog_pol[29]
  PIN gpio_analog_pol[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 775.740 3168.630 776.090 ;
    END
  END gpio_analog_pol[2]
  PIN gpio_analog_pol[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2675.540 0.300 2675.890 ;
    END
  END gpio_analog_pol[30]
  PIN gpio_analog_pol[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2459.540 0.300 2459.890 ;
    END
  END gpio_analog_pol[31]
  PIN gpio_analog_pol[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1821.540 0.300 1821.890 ;
    END
  END gpio_analog_pol[32]
  PIN gpio_analog_pol[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1605.540 0.300 1605.890 ;
    END
  END gpio_analog_pol[33]
  PIN gpio_analog_pol[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1389.540 0.300 1389.890 ;
    END
  END gpio_analog_pol[34]
  PIN gpio_analog_pol[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1173.540 0.300 1173.890 ;
    END
  END gpio_analog_pol[35]
  PIN gpio_analog_pol[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 957.540 0.300 957.890 ;
    END
  END gpio_analog_pol[36]
  PIN gpio_analog_pol[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 741.540 0.300 741.890 ;
    END
  END gpio_analog_pol[37]
  PIN gpio_analog_pol[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.770 -2.000 757.050 0.280 ;
    END
  END gpio_analog_pol[38]
  PIN gpio_analog_pol[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.770 -2.000 1300.050 0.280 ;
    END
  END gpio_analog_pol[39]
  PIN gpio_analog_pol[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1001.740 3168.630 1002.090 ;
    END
  END gpio_analog_pol[3]
  PIN gpio_analog_pol[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.770 -2.000 1574.050 0.280 ;
    END
  END gpio_analog_pol[40]
  PIN gpio_analog_pol[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.770 -2.000 1848.050 0.280 ;
    END
  END gpio_analog_pol[41]
  PIN gpio_analog_pol[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.770 -2.000 2122.050 0.280 ;
    END
  END gpio_analog_pol[42]
  PIN gpio_analog_pol[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 -2.000 2396.050 0.280 ;
    END
  END gpio_analog_pol[43]
  PIN gpio_analog_pol[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1226.740 3168.630 1227.090 ;
    END
  END gpio_analog_pol[4]
  PIN gpio_analog_pol[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1451.740 3168.630 1452.090 ;
    END
  END gpio_analog_pol[5]
  PIN gpio_analog_pol[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1677.740 3168.630 1678.090 ;
    END
  END gpio_analog_pol[6]
  PIN gpio_analog_pol[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2563.740 3168.630 2564.090 ;
    END
  END gpio_analog_pol[7]
  PIN gpio_analog_pol[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2789.740 3168.630 2790.090 ;
    END
  END gpio_analog_pol[8]
  PIN gpio_analog_pol[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3014.740 3168.630 3015.090 ;
    END
  END gpio_analog_pol[9]
  PIN gpio_analog_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 339.920 3168.630 340.270 ;
    END
  END gpio_analog_sel[0]
  PIN gpio_analog_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3255.920 3168.630 3256.270 ;
    END
  END gpio_analog_sel[10]
  PIN gpio_analog_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3480.920 3168.630 3481.270 ;
    END
  END gpio_analog_sel[11]
  PIN gpio_analog_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3705.920 3168.630 3706.270 ;
    END
  END gpio_analog_sel[12]
  PIN gpio_analog_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4151.920 3168.630 4152.270 ;
    END
  END gpio_analog_sel[13]
  PIN gpio_analog_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4597.920 3168.630 4598.270 ;
    END
  END gpio_analog_sel[14]
  PIN gpio_analog_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2948.400 4766.350 2948.680 4768.630 ;
    END
  END gpio_analog_sel[15]
  PIN gpio_analog_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.400 4766.350 2439.680 4768.630 ;
    END
  END gpio_analog_sel[16]
  PIN gpio_analog_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2182.400 4766.350 2182.680 4768.630 ;
    END
  END gpio_analog_sel[17]
  PIN gpio_analog_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.400 4766.350 1737.680 4768.630 ;
    END
  END gpio_analog_sel[18]
  PIN gpio_analog_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.400 4766.350 1228.680 4768.630 ;
    END
  END gpio_analog_sel[19]
  PIN gpio_analog_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 565.920 3168.630 566.270 ;
    END
  END gpio_analog_sel[1]
  PIN gpio_analog_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.400 4766.350 970.680 4768.630 ;
    END
  END gpio_analog_sel[20]
  PIN gpio_analog_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.400 4766.350 713.680 4768.630 ;
    END
  END gpio_analog_sel[21]
  PIN gpio_analog_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.400 4766.350 456.680 4768.630 ;
    END
  END gpio_analog_sel[22]
  PIN gpio_analog_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.400 4766.350 199.680 4768.630 ;
    END
  END gpio_analog_sel[23]
  PIN gpio_analog_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4589.360 0.300 4589.710 ;
    END
  END gpio_analog_sel[24]
  PIN gpio_analog_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3740.360 0.300 3740.710 ;
    END
  END gpio_analog_sel[25]
  PIN gpio_analog_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3524.360 0.300 3524.710 ;
    END
  END gpio_analog_sel[26]
  PIN gpio_analog_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3308.360 0.300 3308.710 ;
    END
  END gpio_analog_sel[27]
  PIN gpio_analog_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3092.360 0.300 3092.710 ;
    END
  END gpio_analog_sel[28]
  PIN gpio_analog_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2876.360 0.300 2876.710 ;
    END
  END gpio_analog_sel[29]
  PIN gpio_analog_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 790.920 3168.630 791.270 ;
    END
  END gpio_analog_sel[2]
  PIN gpio_analog_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2660.360 0.300 2660.710 ;
    END
  END gpio_analog_sel[30]
  PIN gpio_analog_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2444.360 0.300 2444.710 ;
    END
  END gpio_analog_sel[31]
  PIN gpio_analog_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1806.360 0.300 1806.710 ;
    END
  END gpio_analog_sel[32]
  PIN gpio_analog_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1590.360 0.300 1590.710 ;
    END
  END gpio_analog_sel[33]
  PIN gpio_analog_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1374.360 0.300 1374.710 ;
    END
  END gpio_analog_sel[34]
  PIN gpio_analog_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1158.360 0.300 1158.710 ;
    END
  END gpio_analog_sel[35]
  PIN gpio_analog_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 942.360 0.300 942.710 ;
    END
  END gpio_analog_sel[36]
  PIN gpio_analog_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 726.360 0.300 726.710 ;
    END
  END gpio_analog_sel[37]
  PIN gpio_analog_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.950 -2.000 772.230 0.280 ;
    END
  END gpio_analog_sel[38]
  PIN gpio_analog_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.950 -2.000 1315.230 0.280 ;
    END
  END gpio_analog_sel[39]
  PIN gpio_analog_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1016.920 3168.630 1017.270 ;
    END
  END gpio_analog_sel[3]
  PIN gpio_analog_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.950 -2.000 1589.230 0.280 ;
    END
  END gpio_analog_sel[40]
  PIN gpio_analog_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.950 -2.000 1863.230 0.280 ;
    END
  END gpio_analog_sel[41]
  PIN gpio_analog_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.950 -2.000 2137.230 0.280 ;
    END
  END gpio_analog_sel[42]
  PIN gpio_analog_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.950 -2.000 2411.230 0.280 ;
    END
  END gpio_analog_sel[43]
  PIN gpio_analog_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1241.920 3168.630 1242.270 ;
    END
  END gpio_analog_sel[4]
  PIN gpio_analog_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1466.920 3168.630 1467.270 ;
    END
  END gpio_analog_sel[5]
  PIN gpio_analog_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1692.920 3168.630 1693.270 ;
    END
  END gpio_analog_sel[6]
  PIN gpio_analog_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2578.920 3168.630 2579.270 ;
    END
  END gpio_analog_sel[7]
  PIN gpio_analog_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2804.920 3168.630 2805.270 ;
    END
  END gpio_analog_sel[8]
  PIN gpio_analog_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3029.920 3168.630 3030.270 ;
    END
  END gpio_analog_sel[9]
  PIN gpio_dm0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 321.520 3168.630 321.870 ;
    END
  END gpio_dm0[0]
  PIN gpio_dm0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3237.520 3168.630 3237.870 ;
    END
  END gpio_dm0[10]
  PIN gpio_dm0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3462.520 3168.630 3462.870 ;
    END
  END gpio_dm0[11]
  PIN gpio_dm0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3687.520 3168.630 3687.870 ;
    END
  END gpio_dm0[12]
  PIN gpio_dm0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4133.520 3168.630 4133.870 ;
    END
  END gpio_dm0[13]
  PIN gpio_dm0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4579.520 3168.630 4579.870 ;
    END
  END gpio_dm0[14]
  PIN gpio_dm0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2966.800 4766.350 2967.080 4768.630 ;
    END
  END gpio_dm0[15]
  PIN gpio_dm0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2457.800 4766.350 2458.080 4768.630 ;
    END
  END gpio_dm0[16]
  PIN gpio_dm0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2200.800 4766.350 2201.080 4768.630 ;
    END
  END gpio_dm0[17]
  PIN gpio_dm0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.800 4766.350 1756.080 4768.630 ;
    END
  END gpio_dm0[18]
  PIN gpio_dm0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.800 4766.350 1247.080 4768.630 ;
    END
  END gpio_dm0[19]
  PIN gpio_dm0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 547.520 3168.630 547.870 ;
    END
  END gpio_dm0[1]
  PIN gpio_dm0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.800 4766.350 989.080 4768.630 ;
    END
  END gpio_dm0[20]
  PIN gpio_dm0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.800 4766.350 732.080 4768.630 ;
    END
  END gpio_dm0[21]
  PIN gpio_dm0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.800 4766.350 475.080 4768.630 ;
    END
  END gpio_dm0[22]
  PIN gpio_dm0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.800 4766.350 218.080 4768.630 ;
    END
  END gpio_dm0[23]
  PIN gpio_dm0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4607.760 0.300 4608.110 ;
    END
  END gpio_dm0[24]
  PIN gpio_dm0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3758.760 0.300 3759.110 ;
    END
  END gpio_dm0[25]
  PIN gpio_dm0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3542.760 0.300 3543.110 ;
    END
  END gpio_dm0[26]
  PIN gpio_dm0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3326.760 0.300 3327.110 ;
    END
  END gpio_dm0[27]
  PIN gpio_dm0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3110.760 0.300 3111.110 ;
    END
  END gpio_dm0[28]
  PIN gpio_dm0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2894.760 0.300 2895.110 ;
    END
  END gpio_dm0[29]
  PIN gpio_dm0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 772.520 3168.630 772.870 ;
    END
  END gpio_dm0[2]
  PIN gpio_dm0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2678.760 0.300 2679.110 ;
    END
  END gpio_dm0[30]
  PIN gpio_dm0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2462.760 0.300 2463.110 ;
    END
  END gpio_dm0[31]
  PIN gpio_dm0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1824.760 0.300 1825.110 ;
    END
  END gpio_dm0[32]
  PIN gpio_dm0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1608.760 0.300 1609.110 ;
    END
  END gpio_dm0[33]
  PIN gpio_dm0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1392.760 0.300 1393.110 ;
    END
  END gpio_dm0[34]
  PIN gpio_dm0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1176.760 0.300 1177.110 ;
    END
  END gpio_dm0[35]
  PIN gpio_dm0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 960.760 0.300 961.110 ;
    END
  END gpio_dm0[36]
  PIN gpio_dm0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 744.760 0.300 745.110 ;
    END
  END gpio_dm0[37]
  PIN gpio_dm0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.550 -2.000 753.830 0.280 ;
    END
  END gpio_dm0[38]
  PIN gpio_dm0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.550 -2.000 1296.830 0.280 ;
    END
  END gpio_dm0[39]
  PIN gpio_dm0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 998.520 3168.630 998.870 ;
    END
  END gpio_dm0[3]
  PIN gpio_dm0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.550 -2.000 1570.830 0.280 ;
    END
  END gpio_dm0[40]
  PIN gpio_dm0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.550 -2.000 1844.830 0.280 ;
    END
  END gpio_dm0[41]
  PIN gpio_dm0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.550 -2.000 2118.830 0.280 ;
    END
  END gpio_dm0[42]
  PIN gpio_dm0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 -2.000 2392.830 0.280 ;
    END
  END gpio_dm0[43]
  PIN gpio_dm0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1223.520 3168.630 1223.870 ;
    END
  END gpio_dm0[4]
  PIN gpio_dm0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1448.520 3168.630 1448.870 ;
    END
  END gpio_dm0[5]
  PIN gpio_dm0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1674.520 3168.630 1674.870 ;
    END
  END gpio_dm0[6]
  PIN gpio_dm0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2560.520 3168.630 2560.870 ;
    END
  END gpio_dm0[7]
  PIN gpio_dm0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2786.520 3168.630 2786.870 ;
    END
  END gpio_dm0[8]
  PIN gpio_dm0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3011.520 3168.630 3011.870 ;
    END
  END gpio_dm0[9]
  PIN gpio_dm1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 312.320 3168.630 312.670 ;
    END
  END gpio_dm1[0]
  PIN gpio_dm1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3228.320 3168.630 3228.670 ;
    END
  END gpio_dm1[10]
  PIN gpio_dm1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3453.320 3168.630 3453.670 ;
    END
  END gpio_dm1[11]
  PIN gpio_dm1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3678.320 3168.630 3678.670 ;
    END
  END gpio_dm1[12]
  PIN gpio_dm1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4124.320 3168.630 4124.670 ;
    END
  END gpio_dm1[13]
  PIN gpio_dm1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4570.320 3168.630 4570.670 ;
    END
  END gpio_dm1[14]
  PIN gpio_dm1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2976.000 4766.350 2976.280 4768.630 ;
    END
  END gpio_dm1[15]
  PIN gpio_dm1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.000 4766.350 2467.280 4768.630 ;
    END
  END gpio_dm1[16]
  PIN gpio_dm1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.000 4766.350 2210.280 4768.630 ;
    END
  END gpio_dm1[17]
  PIN gpio_dm1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.000 4766.350 1765.280 4768.630 ;
    END
  END gpio_dm1[18]
  PIN gpio_dm1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.000 4766.350 1256.280 4768.630 ;
    END
  END gpio_dm1[19]
  PIN gpio_dm1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 538.320 3168.630 538.670 ;
    END
  END gpio_dm1[1]
  PIN gpio_dm1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.000 4766.350 998.280 4768.630 ;
    END
  END gpio_dm1[20]
  PIN gpio_dm1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.000 4766.350 741.280 4768.630 ;
    END
  END gpio_dm1[21]
  PIN gpio_dm1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.000 4766.350 484.280 4768.630 ;
    END
  END gpio_dm1[22]
  PIN gpio_dm1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.000 4766.350 227.280 4768.630 ;
    END
  END gpio_dm1[23]
  PIN gpio_dm1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4616.960 0.300 4617.310 ;
    END
  END gpio_dm1[24]
  PIN gpio_dm1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3767.960 0.300 3768.310 ;
    END
  END gpio_dm1[25]
  PIN gpio_dm1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3551.960 0.300 3552.310 ;
    END
  END gpio_dm1[26]
  PIN gpio_dm1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3335.960 0.300 3336.310 ;
    END
  END gpio_dm1[27]
  PIN gpio_dm1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3119.960 0.300 3120.310 ;
    END
  END gpio_dm1[28]
  PIN gpio_dm1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2903.960 0.300 2904.310 ;
    END
  END gpio_dm1[29]
  PIN gpio_dm1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 763.320 3168.630 763.670 ;
    END
  END gpio_dm1[2]
  PIN gpio_dm1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2687.960 0.300 2688.310 ;
    END
  END gpio_dm1[30]
  PIN gpio_dm1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2471.960 0.300 2472.310 ;
    END
  END gpio_dm1[31]
  PIN gpio_dm1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1833.960 0.300 1834.310 ;
    END
  END gpio_dm1[32]
  PIN gpio_dm1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1617.960 0.300 1618.310 ;
    END
  END gpio_dm1[33]
  PIN gpio_dm1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1401.960 0.300 1402.310 ;
    END
  END gpio_dm1[34]
  PIN gpio_dm1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1185.960 0.300 1186.310 ;
    END
  END gpio_dm1[35]
  PIN gpio_dm1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 969.960 0.300 970.310 ;
    END
  END gpio_dm1[36]
  PIN gpio_dm1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 753.960 0.300 754.310 ;
    END
  END gpio_dm1[37]
  PIN gpio_dm1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.350 -2.000 744.630 0.280 ;
    END
  END gpio_dm1[38]
  PIN gpio_dm1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.350 -2.000 1287.630 0.280 ;
    END
  END gpio_dm1[39]
  PIN gpio_dm1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 989.320 3168.630 989.670 ;
    END
  END gpio_dm1[3]
  PIN gpio_dm1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.350 -2.000 1561.630 0.280 ;
    END
  END gpio_dm1[40]
  PIN gpio_dm1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.350 -2.000 1835.630 0.280 ;
    END
  END gpio_dm1[41]
  PIN gpio_dm1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.350 -2.000 2109.630 0.280 ;
    END
  END gpio_dm1[42]
  PIN gpio_dm1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2383.350 -2.000 2383.630 0.280 ;
    END
  END gpio_dm1[43]
  PIN gpio_dm1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1214.320 3168.630 1214.670 ;
    END
  END gpio_dm1[4]
  PIN gpio_dm1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1439.320 3168.630 1439.670 ;
    END
  END gpio_dm1[5]
  PIN gpio_dm1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1665.320 3168.630 1665.670 ;
    END
  END gpio_dm1[6]
  PIN gpio_dm1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2551.320 3168.630 2551.670 ;
    END
  END gpio_dm1[7]
  PIN gpio_dm1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2777.320 3168.630 2777.670 ;
    END
  END gpio_dm1[8]
  PIN gpio_dm1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3002.320 3168.630 3002.670 ;
    END
  END gpio_dm1[9]
  PIN gpio_dm2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 343.140 3168.630 343.490 ;
    END
  END gpio_dm2[0]
  PIN gpio_dm2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3259.140 3168.630 3259.490 ;
    END
  END gpio_dm2[10]
  PIN gpio_dm2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3484.140 3168.630 3484.490 ;
    END
  END gpio_dm2[11]
  PIN gpio_dm2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3709.140 3168.630 3709.490 ;
    END
  END gpio_dm2[12]
  PIN gpio_dm2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4155.140 3168.630 4155.490 ;
    END
  END gpio_dm2[13]
  PIN gpio_dm2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4601.140 3168.630 4601.490 ;
    END
  END gpio_dm2[14]
  PIN gpio_dm2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2945.180 4766.350 2945.460 4768.630 ;
    END
  END gpio_dm2[15]
  PIN gpio_dm2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2436.180 4766.350 2436.460 4768.630 ;
    END
  END gpio_dm2[16]
  PIN gpio_dm2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.180 4766.350 2179.460 4768.630 ;
    END
  END gpio_dm2[17]
  PIN gpio_dm2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.180 4766.350 1734.460 4768.630 ;
    END
  END gpio_dm2[18]
  PIN gpio_dm2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.180 4766.350 1225.460 4768.630 ;
    END
  END gpio_dm2[19]
  PIN gpio_dm2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 569.140 3168.630 569.490 ;
    END
  END gpio_dm2[1]
  PIN gpio_dm2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.180 4766.350 967.460 4768.630 ;
    END
  END gpio_dm2[20]
  PIN gpio_dm2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.180 4766.350 710.460 4768.630 ;
    END
  END gpio_dm2[21]
  PIN gpio_dm2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.180 4766.350 453.460 4768.630 ;
    END
  END gpio_dm2[22]
  PIN gpio_dm2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.180 4766.350 196.460 4768.630 ;
    END
  END gpio_dm2[23]
  PIN gpio_dm2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4586.140 0.300 4586.490 ;
    END
  END gpio_dm2[24]
  PIN gpio_dm2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3737.140 0.300 3737.490 ;
    END
  END gpio_dm2[25]
  PIN gpio_dm2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3521.140 0.300 3521.490 ;
    END
  END gpio_dm2[26]
  PIN gpio_dm2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3305.140 0.300 3305.490 ;
    END
  END gpio_dm2[27]
  PIN gpio_dm2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3089.140 0.300 3089.490 ;
    END
  END gpio_dm2[28]
  PIN gpio_dm2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2873.140 0.300 2873.490 ;
    END
  END gpio_dm2[29]
  PIN gpio_dm2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 794.140 3168.630 794.490 ;
    END
  END gpio_dm2[2]
  PIN gpio_dm2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2657.140 0.300 2657.490 ;
    END
  END gpio_dm2[30]
  PIN gpio_dm2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2441.140 0.300 2441.490 ;
    END
  END gpio_dm2[31]
  PIN gpio_dm2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1803.140 0.300 1803.490 ;
    END
  END gpio_dm2[32]
  PIN gpio_dm2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1587.140 0.300 1587.490 ;
    END
  END gpio_dm2[33]
  PIN gpio_dm2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1371.140 0.300 1371.490 ;
    END
  END gpio_dm2[34]
  PIN gpio_dm2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1155.140 0.300 1155.490 ;
    END
  END gpio_dm2[35]
  PIN gpio_dm2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 939.140 0.300 939.490 ;
    END
  END gpio_dm2[36]
  PIN gpio_dm2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 723.140 0.300 723.490 ;
    END
  END gpio_dm2[37]
  PIN gpio_dm2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.170 -2.000 775.450 0.280 ;
    END
  END gpio_dm2[38]
  PIN gpio_dm2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.170 -2.000 1318.450 0.280 ;
    END
  END gpio_dm2[39]
  PIN gpio_dm2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1020.140 3168.630 1020.490 ;
    END
  END gpio_dm2[3]
  PIN gpio_dm2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.170 -2.000 1592.450 0.280 ;
    END
  END gpio_dm2[40]
  PIN gpio_dm2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.170 -2.000 1866.450 0.280 ;
    END
  END gpio_dm2[41]
  PIN gpio_dm2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.170 -2.000 2140.450 0.280 ;
    END
  END gpio_dm2[42]
  PIN gpio_dm2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.170 -2.000 2414.450 0.280 ;
    END
  END gpio_dm2[43]
  PIN gpio_dm2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1245.140 3168.630 1245.490 ;
    END
  END gpio_dm2[4]
  PIN gpio_dm2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1470.140 3168.630 1470.490 ;
    END
  END gpio_dm2[5]
  PIN gpio_dm2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1696.140 3168.630 1696.490 ;
    END
  END gpio_dm2[6]
  PIN gpio_dm2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2582.140 3168.630 2582.490 ;
    END
  END gpio_dm2[7]
  PIN gpio_dm2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2808.140 3168.630 2808.490 ;
    END
  END gpio_dm2[8]
  PIN gpio_dm2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3033.140 3168.630 3033.490 ;
    END
  END gpio_dm2[9]
  PIN gpio_holdover[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 346.360 3168.630 346.710 ;
    END
  END gpio_holdover[0]
  PIN gpio_holdover[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3262.360 3168.630 3262.710 ;
    END
  END gpio_holdover[10]
  PIN gpio_holdover[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3487.360 3168.630 3487.710 ;
    END
  END gpio_holdover[11]
  PIN gpio_holdover[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3712.360 3168.630 3712.710 ;
    END
  END gpio_holdover[12]
  PIN gpio_holdover[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4158.360 3168.630 4158.710 ;
    END
  END gpio_holdover[13]
  PIN gpio_holdover[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4604.360 3168.630 4604.710 ;
    END
  END gpio_holdover[14]
  PIN gpio_holdover[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2941.960 4766.350 2942.240 4768.630 ;
    END
  END gpio_holdover[15]
  PIN gpio_holdover[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2432.960 4766.350 2433.240 4768.630 ;
    END
  END gpio_holdover[16]
  PIN gpio_holdover[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.960 4766.350 2176.240 4768.630 ;
    END
  END gpio_holdover[17]
  PIN gpio_holdover[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.960 4766.350 1731.240 4768.630 ;
    END
  END gpio_holdover[18]
  PIN gpio_holdover[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.960 4766.350 1222.240 4768.630 ;
    END
  END gpio_holdover[19]
  PIN gpio_holdover[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 572.360 3168.630 572.710 ;
    END
  END gpio_holdover[1]
  PIN gpio_holdover[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.960 4766.350 964.240 4768.630 ;
    END
  END gpio_holdover[20]
  PIN gpio_holdover[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.960 4766.350 707.240 4768.630 ;
    END
  END gpio_holdover[21]
  PIN gpio_holdover[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.960 4766.350 450.240 4768.630 ;
    END
  END gpio_holdover[22]
  PIN gpio_holdover[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.960 4766.350 193.240 4768.630 ;
    END
  END gpio_holdover[23]
  PIN gpio_holdover[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4582.920 0.300 4583.270 ;
    END
  END gpio_holdover[24]
  PIN gpio_holdover[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3733.920 0.300 3734.270 ;
    END
  END gpio_holdover[25]
  PIN gpio_holdover[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3517.920 0.300 3518.270 ;
    END
  END gpio_holdover[26]
  PIN gpio_holdover[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3301.920 0.300 3302.270 ;
    END
  END gpio_holdover[27]
  PIN gpio_holdover[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3085.920 0.300 3086.270 ;
    END
  END gpio_holdover[28]
  PIN gpio_holdover[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2869.920 0.300 2870.270 ;
    END
  END gpio_holdover[29]
  PIN gpio_holdover[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 797.360 3168.630 797.710 ;
    END
  END gpio_holdover[2]
  PIN gpio_holdover[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2653.920 0.300 2654.270 ;
    END
  END gpio_holdover[30]
  PIN gpio_holdover[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2437.920 0.300 2438.270 ;
    END
  END gpio_holdover[31]
  PIN gpio_holdover[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1799.920 0.300 1800.270 ;
    END
  END gpio_holdover[32]
  PIN gpio_holdover[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1583.920 0.300 1584.270 ;
    END
  END gpio_holdover[33]
  PIN gpio_holdover[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1367.920 0.300 1368.270 ;
    END
  END gpio_holdover[34]
  PIN gpio_holdover[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1151.920 0.300 1152.270 ;
    END
  END gpio_holdover[35]
  PIN gpio_holdover[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 935.920 0.300 936.270 ;
    END
  END gpio_holdover[36]
  PIN gpio_holdover[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 719.920 0.300 720.270 ;
    END
  END gpio_holdover[37]
  PIN gpio_holdover[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.390 -2.000 778.670 0.280 ;
    END
  END gpio_holdover[38]
  PIN gpio_holdover[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.390 -2.000 1321.670 0.280 ;
    END
  END gpio_holdover[39]
  PIN gpio_holdover[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1023.360 3168.630 1023.710 ;
    END
  END gpio_holdover[3]
  PIN gpio_holdover[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.390 -2.000 1595.670 0.280 ;
    END
  END gpio_holdover[40]
  PIN gpio_holdover[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.390 -2.000 1869.670 0.280 ;
    END
  END gpio_holdover[41]
  PIN gpio_holdover[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.390 -2.000 2143.670 0.280 ;
    END
  END gpio_holdover[42]
  PIN gpio_holdover[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.390 -2.000 2417.670 0.280 ;
    END
  END gpio_holdover[43]
  PIN gpio_holdover[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1248.360 3168.630 1248.710 ;
    END
  END gpio_holdover[4]
  PIN gpio_holdover[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1473.360 3168.630 1473.710 ;
    END
  END gpio_holdover[5]
  PIN gpio_holdover[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1699.360 3168.630 1699.710 ;
    END
  END gpio_holdover[6]
  PIN gpio_holdover[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2585.360 3168.630 2585.710 ;
    END
  END gpio_holdover[7]
  PIN gpio_holdover[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2811.360 3168.630 2811.710 ;
    END
  END gpio_holdover[8]
  PIN gpio_holdover[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3036.360 3168.630 3036.710 ;
    END
  END gpio_holdover[9]
  PIN gpio_ib_mode_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 361.540 3168.630 361.890 ;
    END
  END gpio_ib_mode_sel[0]
  PIN gpio_ib_mode_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3277.540 3168.630 3277.890 ;
    END
  END gpio_ib_mode_sel[10]
  PIN gpio_ib_mode_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3502.540 3168.630 3502.890 ;
    END
  END gpio_ib_mode_sel[11]
  PIN gpio_ib_mode_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3727.540 3168.630 3727.890 ;
    END
  END gpio_ib_mode_sel[12]
  PIN gpio_ib_mode_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4173.540 3168.630 4173.890 ;
    END
  END gpio_ib_mode_sel[13]
  PIN gpio_ib_mode_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4619.540 3168.630 4619.890 ;
    END
  END gpio_ib_mode_sel[14]
  PIN gpio_ib_mode_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2926.780 4766.350 2927.060 4768.630 ;
    END
  END gpio_ib_mode_sel[15]
  PIN gpio_ib_mode_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.780 4766.350 2418.060 4768.630 ;
    END
  END gpio_ib_mode_sel[16]
  PIN gpio_ib_mode_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.780 4766.350 2161.060 4768.630 ;
    END
  END gpio_ib_mode_sel[17]
  PIN gpio_ib_mode_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.780 4766.350 1716.060 4768.630 ;
    END
  END gpio_ib_mode_sel[18]
  PIN gpio_ib_mode_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.780 4766.350 1207.060 4768.630 ;
    END
  END gpio_ib_mode_sel[19]
  PIN gpio_ib_mode_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 587.540 3168.630 587.890 ;
    END
  END gpio_ib_mode_sel[1]
  PIN gpio_ib_mode_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.780 4766.350 949.060 4768.630 ;
    END
  END gpio_ib_mode_sel[20]
  PIN gpio_ib_mode_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.780 4766.350 692.060 4768.630 ;
    END
  END gpio_ib_mode_sel[21]
  PIN gpio_ib_mode_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.780 4766.350 435.060 4768.630 ;
    END
  END gpio_ib_mode_sel[22]
  PIN gpio_ib_mode_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.780 4766.350 178.060 4768.630 ;
    END
  END gpio_ib_mode_sel[23]
  PIN gpio_ib_mode_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4567.740 0.300 4568.090 ;
    END
  END gpio_ib_mode_sel[24]
  PIN gpio_ib_mode_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3718.740 0.300 3719.090 ;
    END
  END gpio_ib_mode_sel[25]
  PIN gpio_ib_mode_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3502.740 0.300 3503.090 ;
    END
  END gpio_ib_mode_sel[26]
  PIN gpio_ib_mode_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3286.740 0.300 3287.090 ;
    END
  END gpio_ib_mode_sel[27]
  PIN gpio_ib_mode_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3070.740 0.300 3071.090 ;
    END
  END gpio_ib_mode_sel[28]
  PIN gpio_ib_mode_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2854.740 0.300 2855.090 ;
    END
  END gpio_ib_mode_sel[29]
  PIN gpio_ib_mode_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 812.540 3168.630 812.890 ;
    END
  END gpio_ib_mode_sel[2]
  PIN gpio_ib_mode_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2638.740 0.300 2639.090 ;
    END
  END gpio_ib_mode_sel[30]
  PIN gpio_ib_mode_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2422.740 0.300 2423.090 ;
    END
  END gpio_ib_mode_sel[31]
  PIN gpio_ib_mode_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1784.740 0.300 1785.090 ;
    END
  END gpio_ib_mode_sel[32]
  PIN gpio_ib_mode_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1568.740 0.300 1569.090 ;
    END
  END gpio_ib_mode_sel[33]
  PIN gpio_ib_mode_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1352.740 0.300 1353.090 ;
    END
  END gpio_ib_mode_sel[34]
  PIN gpio_ib_mode_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1136.740 0.300 1137.090 ;
    END
  END gpio_ib_mode_sel[35]
  PIN gpio_ib_mode_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 920.740 0.300 921.090 ;
    END
  END gpio_ib_mode_sel[36]
  PIN gpio_ib_mode_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 704.740 0.300 705.090 ;
    END
  END gpio_ib_mode_sel[37]
  PIN gpio_ib_mode_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.570 -2.000 793.850 0.280 ;
    END
  END gpio_ib_mode_sel[38]
  PIN gpio_ib_mode_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.570 -2.000 1336.850 0.280 ;
    END
  END gpio_ib_mode_sel[39]
  PIN gpio_ib_mode_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1038.540 3168.630 1038.890 ;
    END
  END gpio_ib_mode_sel[3]
  PIN gpio_ib_mode_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.570 -2.000 1610.850 0.280 ;
    END
  END gpio_ib_mode_sel[40]
  PIN gpio_ib_mode_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1884.570 -2.000 1884.850 0.280 ;
    END
  END gpio_ib_mode_sel[41]
  PIN gpio_ib_mode_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.570 -2.000 2158.850 0.280 ;
    END
  END gpio_ib_mode_sel[42]
  PIN gpio_ib_mode_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2432.570 -2.000 2432.850 0.280 ;
    END
  END gpio_ib_mode_sel[43]
  PIN gpio_ib_mode_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1263.540 3168.630 1263.890 ;
    END
  END gpio_ib_mode_sel[4]
  PIN gpio_ib_mode_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1488.540 3168.630 1488.890 ;
    END
  END gpio_ib_mode_sel[5]
  PIN gpio_ib_mode_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1714.540 3168.630 1714.890 ;
    END
  END gpio_ib_mode_sel[6]
  PIN gpio_ib_mode_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2600.540 3168.630 2600.890 ;
    END
  END gpio_ib_mode_sel[7]
  PIN gpio_ib_mode_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2826.540 3168.630 2826.890 ;
    END
  END gpio_ib_mode_sel[8]
  PIN gpio_ib_mode_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3051.540 3168.630 3051.890 ;
    END
  END gpio_ib_mode_sel[9]
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 293.920 3168.630 294.270 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3209.920 3168.630 3210.270 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3434.920 3168.630 3435.270 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3659.920 3168.630 3660.270 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4105.920 3168.630 4106.270 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4551.920 3168.630 4552.270 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2994.400 4766.350 2994.680 4768.630 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.400 4766.350 2485.680 4768.630 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.400 4766.350 2228.680 4768.630 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.400 4766.350 1783.680 4768.630 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.400 4766.350 1274.680 4768.630 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 519.920 3168.630 520.270 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.400 4766.350 1016.680 4768.630 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.400 4766.350 759.680 4768.630 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.400 4766.350 502.680 4768.630 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.400 4766.350 245.680 4768.630 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4635.360 0.300 4635.710 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3786.360 0.300 3786.710 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3570.360 0.300 3570.710 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3354.360 0.300 3354.710 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3138.360 0.300 3138.710 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2922.360 0.300 2922.710 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 744.920 3168.630 745.270 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2706.360 0.300 2706.710 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2490.360 0.300 2490.710 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1852.360 0.300 1852.710 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1636.360 0.300 1636.710 ;
    END
  END gpio_in[33]
  PIN gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1420.360 0.300 1420.710 ;
    END
  END gpio_in[34]
  PIN gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1204.360 0.300 1204.710 ;
    END
  END gpio_in[35]
  PIN gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 988.360 0.300 988.710 ;
    END
  END gpio_in[36]
  PIN gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 772.360 0.300 772.710 ;
    END
  END gpio_in[37]
  PIN gpio_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.950 -2.000 726.230 0.280 ;
    END
  END gpio_in[38]
  PIN gpio_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.950 -2.000 1269.230 0.280 ;
    END
  END gpio_in[39]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 970.920 3168.630 971.270 ;
    END
  END gpio_in[3]
  PIN gpio_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.950 -2.000 1543.230 0.280 ;
    END
  END gpio_in[40]
  PIN gpio_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.950 -2.000 1817.230 0.280 ;
    END
  END gpio_in[41]
  PIN gpio_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.950 -2.000 2091.230 0.280 ;
    END
  END gpio_in[42]
  PIN gpio_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.950 -2.000 2365.230 0.280 ;
    END
  END gpio_in[43]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1195.920 3168.630 1196.270 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1420.920 3168.630 1421.270 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1646.920 3168.630 1647.270 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2532.920 3168.630 2533.270 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2758.920 3168.630 2759.270 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2983.920 3168.630 2984.270 ;
    END
  END gpio_in[9]
  PIN gpio_in_h[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 367.520 3168.630 367.870 ;
    END
  END gpio_in_h[0]
  PIN gpio_in_h[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3283.520 3168.630 3283.870 ;
    END
  END gpio_in_h[10]
  PIN gpio_in_h[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3508.520 3168.630 3508.870 ;
    END
  END gpio_in_h[11]
  PIN gpio_in_h[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3733.520 3168.630 3733.870 ;
    END
  END gpio_in_h[12]
  PIN gpio_in_h[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4179.520 3168.630 4179.870 ;
    END
  END gpio_in_h[13]
  PIN gpio_in_h[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4625.520 3168.630 4625.870 ;
    END
  END gpio_in_h[14]
  PIN gpio_in_h[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2920.800 4766.350 2921.080 4768.630 ;
    END
  END gpio_in_h[15]
  PIN gpio_in_h[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.800 4766.350 2412.080 4768.630 ;
    END
  END gpio_in_h[16]
  PIN gpio_in_h[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.800 4766.350 2155.080 4768.630 ;
    END
  END gpio_in_h[17]
  PIN gpio_in_h[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.800 4766.350 1710.080 4768.630 ;
    END
  END gpio_in_h[18]
  PIN gpio_in_h[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.800 4766.350 1201.080 4768.630 ;
    END
  END gpio_in_h[19]
  PIN gpio_in_h[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 593.520 3168.630 593.870 ;
    END
  END gpio_in_h[1]
  PIN gpio_in_h[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.800 4766.350 943.080 4768.630 ;
    END
  END gpio_in_h[20]
  PIN gpio_in_h[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.800 4766.350 686.080 4768.630 ;
    END
  END gpio_in_h[21]
  PIN gpio_in_h[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.800 4766.350 429.080 4768.630 ;
    END
  END gpio_in_h[22]
  PIN gpio_in_h[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.800 4766.350 172.080 4768.630 ;
    END
  END gpio_in_h[23]
  PIN gpio_in_h[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4561.760 0.300 4562.110 ;
    END
  END gpio_in_h[24]
  PIN gpio_in_h[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3712.760 0.300 3713.110 ;
    END
  END gpio_in_h[25]
  PIN gpio_in_h[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3496.760 0.300 3497.110 ;
    END
  END gpio_in_h[26]
  PIN gpio_in_h[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3280.760 0.300 3281.110 ;
    END
  END gpio_in_h[27]
  PIN gpio_in_h[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3064.760 0.300 3065.110 ;
    END
  END gpio_in_h[28]
  PIN gpio_in_h[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2848.760 0.300 2849.110 ;
    END
  END gpio_in_h[29]
  PIN gpio_in_h[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 818.520 3168.630 818.870 ;
    END
  END gpio_in_h[2]
  PIN gpio_in_h[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2632.760 0.300 2633.110 ;
    END
  END gpio_in_h[30]
  PIN gpio_in_h[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2416.760 0.300 2417.110 ;
    END
  END gpio_in_h[31]
  PIN gpio_in_h[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1778.760 0.300 1779.110 ;
    END
  END gpio_in_h[32]
  PIN gpio_in_h[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1562.760 0.300 1563.110 ;
    END
  END gpio_in_h[33]
  PIN gpio_in_h[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1346.760 0.300 1347.110 ;
    END
  END gpio_in_h[34]
  PIN gpio_in_h[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1130.760 0.300 1131.110 ;
    END
  END gpio_in_h[35]
  PIN gpio_in_h[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 914.760 0.300 915.110 ;
    END
  END gpio_in_h[36]
  PIN gpio_in_h[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 698.760 0.300 699.110 ;
    END
  END gpio_in_h[37]
  PIN gpio_in_h[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.550 -2.000 799.830 0.280 ;
    END
  END gpio_in_h[38]
  PIN gpio_in_h[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.550 -2.000 1342.830 0.280 ;
    END
  END gpio_in_h[39]
  PIN gpio_in_h[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1044.520 3168.630 1044.870 ;
    END
  END gpio_in_h[3]
  PIN gpio_in_h[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.550 -2.000 1616.830 0.280 ;
    END
  END gpio_in_h[40]
  PIN gpio_in_h[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.550 -2.000 1890.830 0.280 ;
    END
  END gpio_in_h[41]
  PIN gpio_in_h[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.550 -2.000 2164.830 0.280 ;
    END
  END gpio_in_h[42]
  PIN gpio_in_h[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2438.550 -2.000 2438.830 0.280 ;
    END
  END gpio_in_h[43]
  PIN gpio_in_h[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1269.520 3168.630 1269.870 ;
    END
  END gpio_in_h[4]
  PIN gpio_in_h[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1494.520 3168.630 1494.870 ;
    END
  END gpio_in_h[5]
  PIN gpio_in_h[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1720.520 3168.630 1720.870 ;
    END
  END gpio_in_h[6]
  PIN gpio_in_h[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2606.520 3168.630 2606.870 ;
    END
  END gpio_in_h[7]
  PIN gpio_in_h[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2832.520 3168.630 2832.870 ;
    END
  END gpio_in_h[8]
  PIN gpio_in_h[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3057.520 3168.630 3057.870 ;
    END
  END gpio_in_h[9]
  PIN gpio_inp_dis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 327.500 3168.630 327.850 ;
    END
  END gpio_inp_dis[0]
  PIN gpio_inp_dis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3243.500 3168.630 3243.850 ;
    END
  END gpio_inp_dis[10]
  PIN gpio_inp_dis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3468.500 3168.630 3468.850 ;
    END
  END gpio_inp_dis[11]
  PIN gpio_inp_dis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3693.500 3168.630 3693.850 ;
    END
  END gpio_inp_dis[12]
  PIN gpio_inp_dis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4139.500 3168.630 4139.850 ;
    END
  END gpio_inp_dis[13]
  PIN gpio_inp_dis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4585.500 3168.630 4585.850 ;
    END
  END gpio_inp_dis[14]
  PIN gpio_inp_dis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2960.820 4766.350 2961.100 4768.630 ;
    END
  END gpio_inp_dis[15]
  PIN gpio_inp_dis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.820 4766.350 2452.100 4768.630 ;
    END
  END gpio_inp_dis[16]
  PIN gpio_inp_dis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.820 4766.350 2195.100 4768.630 ;
    END
  END gpio_inp_dis[17]
  PIN gpio_inp_dis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.820 4766.350 1750.100 4768.630 ;
    END
  END gpio_inp_dis[18]
  PIN gpio_inp_dis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.820 4766.350 1241.100 4768.630 ;
    END
  END gpio_inp_dis[19]
  PIN gpio_inp_dis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 553.500 3168.630 553.850 ;
    END
  END gpio_inp_dis[1]
  PIN gpio_inp_dis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.820 4766.350 983.100 4768.630 ;
    END
  END gpio_inp_dis[20]
  PIN gpio_inp_dis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.820 4766.350 726.100 4768.630 ;
    END
  END gpio_inp_dis[21]
  PIN gpio_inp_dis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.820 4766.350 469.100 4768.630 ;
    END
  END gpio_inp_dis[22]
  PIN gpio_inp_dis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.820 4766.350 212.100 4768.630 ;
    END
  END gpio_inp_dis[23]
  PIN gpio_inp_dis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4601.780 0.300 4602.130 ;
    END
  END gpio_inp_dis[24]
  PIN gpio_inp_dis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3752.780 0.300 3753.130 ;
    END
  END gpio_inp_dis[25]
  PIN gpio_inp_dis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3536.780 0.300 3537.130 ;
    END
  END gpio_inp_dis[26]
  PIN gpio_inp_dis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3320.780 0.300 3321.130 ;
    END
  END gpio_inp_dis[27]
  PIN gpio_inp_dis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3104.780 0.300 3105.130 ;
    END
  END gpio_inp_dis[28]
  PIN gpio_inp_dis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2888.780 0.300 2889.130 ;
    END
  END gpio_inp_dis[29]
  PIN gpio_inp_dis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 778.500 3168.630 778.850 ;
    END
  END gpio_inp_dis[2]
  PIN gpio_inp_dis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2672.780 0.300 2673.130 ;
    END
  END gpio_inp_dis[30]
  PIN gpio_inp_dis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2456.780 0.300 2457.130 ;
    END
  END gpio_inp_dis[31]
  PIN gpio_inp_dis[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1818.780 0.300 1819.130 ;
    END
  END gpio_inp_dis[32]
  PIN gpio_inp_dis[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1602.780 0.300 1603.130 ;
    END
  END gpio_inp_dis[33]
  PIN gpio_inp_dis[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1386.780 0.300 1387.130 ;
    END
  END gpio_inp_dis[34]
  PIN gpio_inp_dis[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1170.780 0.300 1171.130 ;
    END
  END gpio_inp_dis[35]
  PIN gpio_inp_dis[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 954.780 0.300 955.130 ;
    END
  END gpio_inp_dis[36]
  PIN gpio_inp_dis[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 738.780 0.300 739.130 ;
    END
  END gpio_inp_dis[37]
  PIN gpio_inp_dis[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.530 -2.000 759.810 0.280 ;
    END
  END gpio_inp_dis[38]
  PIN gpio_inp_dis[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.530 -2.000 1302.810 0.280 ;
    END
  END gpio_inp_dis[39]
  PIN gpio_inp_dis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1004.500 3168.630 1004.850 ;
    END
  END gpio_inp_dis[3]
  PIN gpio_inp_dis[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.530 -2.000 1576.810 0.280 ;
    END
  END gpio_inp_dis[40]
  PIN gpio_inp_dis[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.530 -2.000 1850.810 0.280 ;
    END
  END gpio_inp_dis[41]
  PIN gpio_inp_dis[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.530 -2.000 2124.810 0.280 ;
    END
  END gpio_inp_dis[42]
  PIN gpio_inp_dis[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.530 -2.000 2398.810 0.280 ;
    END
  END gpio_inp_dis[43]
  PIN gpio_inp_dis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1229.500 3168.630 1229.850 ;
    END
  END gpio_inp_dis[4]
  PIN gpio_inp_dis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1454.500 3168.630 1454.850 ;
    END
  END gpio_inp_dis[5]
  PIN gpio_inp_dis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1680.500 3168.630 1680.850 ;
    END
  END gpio_inp_dis[6]
  PIN gpio_inp_dis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2566.500 3168.630 2566.850 ;
    END
  END gpio_inp_dis[7]
  PIN gpio_inp_dis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2792.500 3168.630 2792.850 ;
    END
  END gpio_inp_dis[8]
  PIN gpio_inp_dis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3017.500 3168.630 3017.850 ;
    END
  END gpio_inp_dis[9]
  PIN gpio_loopback_one[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 380.025 3168.630 380.335 ;
    END
  END gpio_loopback_one[0]
  PIN gpio_loopback_one[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3290.030 3168.630 3290.340 ;
    END
  END gpio_loopback_one[10]
  PIN gpio_loopback_one[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3515.030 3168.630 3515.340 ;
    END
  END gpio_loopback_one[11]
  PIN gpio_loopback_one[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3740.030 3168.630 3740.340 ;
    END
  END gpio_loopback_one[12]
  PIN gpio_loopback_one[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4185.030 3168.630 4185.340 ;
    END
  END gpio_loopback_one[13]
  PIN gpio_loopback_one[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4635.030 3168.630 4635.340 ;
    END
  END gpio_loopback_one[14]
  PIN gpio_loopback_one[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2891.490 4766.350 2891.790 4768.630 ;
    END
  END gpio_loopback_one[15]
  PIN gpio_loopback_one[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2394.490 4766.350 2394.790 4768.630 ;
    END
  END gpio_loopback_one[16]
  PIN gpio_loopback_one[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.490 4766.350 2138.790 4768.630 ;
    END
  END gpio_loopback_one[17]
  PIN gpio_loopback_one[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.490 4766.350 1693.790 4768.630 ;
    END
  END gpio_loopback_one[18]
  PIN gpio_loopback_one[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.490 4766.350 1171.790 4768.630 ;
    END
  END gpio_loopback_one[19]
  PIN gpio_loopback_one[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 605.025 3168.630 605.335 ;
    END
  END gpio_loopback_one[1]
  PIN gpio_loopback_one[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 4766.350 915.790 4768.630 ;
    END
  END gpio_loopback_one[20]
  PIN gpio_loopback_one[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.490 4766.350 659.790 4768.630 ;
    END
  END gpio_loopback_one[21]
  PIN gpio_loopback_one[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.490 4766.350 403.790 4768.630 ;
    END
  END gpio_loopback_one[22]
  PIN gpio_loopback_one[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.490 4766.350 147.790 4768.630 ;
    END
  END gpio_loopback_one[23]
  PIN gpio_loopback_one[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4533.220 0.300 4533.520 ;
    END
  END gpio_loopback_one[24]
  PIN gpio_loopback_one[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3683.220 0.300 3683.520 ;
    END
  END gpio_loopback_one[25]
  PIN gpio_loopback_one[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3468.220 0.300 3468.520 ;
    END
  END gpio_loopback_one[26]
  PIN gpio_loopback_one[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3253.220 0.300 3253.520 ;
    END
  END gpio_loopback_one[27]
  PIN gpio_loopback_one[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3038.220 0.300 3038.520 ;
    END
  END gpio_loopback_one[28]
  PIN gpio_loopback_one[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2823.220 0.300 2823.520 ;
    END
  END gpio_loopback_one[29]
  PIN gpio_loopback_one[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 830.025 3168.630 830.335 ;
    END
  END gpio_loopback_one[2]
  PIN gpio_loopback_one[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2608.220 0.300 2608.520 ;
    END
  END gpio_loopback_one[30]
  PIN gpio_loopback_one[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2393.220 0.300 2393.520 ;
    END
  END gpio_loopback_one[31]
  PIN gpio_loopback_one[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1748.220 0.300 1748.520 ;
    END
  END gpio_loopback_one[32]
  PIN gpio_loopback_one[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1533.220 0.300 1533.520 ;
    END
  END gpio_loopback_one[33]
  PIN gpio_loopback_one[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1318.220 0.300 1318.520 ;
    END
  END gpio_loopback_one[34]
  PIN gpio_loopback_one[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1103.220 0.300 1103.520 ;
    END
  END gpio_loopback_one[35]
  PIN gpio_loopback_one[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 888.220 0.300 888.520 ;
    END
  END gpio_loopback_one[36]
  PIN gpio_loopback_one[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 673.220 0.300 673.520 ;
    END
  END gpio_loopback_one[37]
  PIN gpio_loopback_one[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.900 -2.000 803.160 0.280 ;
    END
  END gpio_loopback_one[38]
  PIN gpio_loopback_one[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.900 -2.000 1346.160 0.280 ;
    END
  END gpio_loopback_one[39]
  PIN gpio_loopback_one[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1055.025 3168.630 1055.335 ;
    END
  END gpio_loopback_one[3]
  PIN gpio_loopback_one[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.900 -2.000 1620.160 0.280 ;
    END
  END gpio_loopback_one[40]
  PIN gpio_loopback_one[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.900 -2.000 1894.160 0.280 ;
    END
  END gpio_loopback_one[41]
  PIN gpio_loopback_one[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.900 -2.000 2168.160 0.280 ;
    END
  END gpio_loopback_one[42]
  PIN gpio_loopback_one[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.900 -2.000 2442.160 0.280 ;
    END
  END gpio_loopback_one[43]
  PIN gpio_loopback_one[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1280.025 3168.630 1280.335 ;
    END
  END gpio_loopback_one[4]
  PIN gpio_loopback_one[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1505.025 3168.630 1505.335 ;
    END
  END gpio_loopback_one[5]
  PIN gpio_loopback_one[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1730.025 3168.630 1730.335 ;
    END
  END gpio_loopback_one[6]
  PIN gpio_loopback_one[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2615.025 3168.630 2615.335 ;
    END
  END gpio_loopback_one[7]
  PIN gpio_loopback_one[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2840.030 3168.630 2840.340 ;
    END
  END gpio_loopback_one[8]
  PIN gpio_loopback_one[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3065.030 3168.630 3065.340 ;
    END
  END gpio_loopback_one[9]
  PIN gpio_loopback_zero[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 390.030 3168.630 390.340 ;
    END
  END gpio_loopback_zero[0]
  PIN gpio_loopback_zero[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3300.030 3168.630 3300.340 ;
    END
  END gpio_loopback_zero[10]
  PIN gpio_loopback_zero[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3525.030 3168.630 3525.340 ;
    END
  END gpio_loopback_zero[11]
  PIN gpio_loopback_zero[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3750.030 3168.630 3750.340 ;
    END
  END gpio_loopback_zero[12]
  PIN gpio_loopback_zero[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4195.030 3168.630 4195.340 ;
    END
  END gpio_loopback_zero[13]
  PIN gpio_loopback_zero[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4645.030 3168.630 4645.340 ;
    END
  END gpio_loopback_zero[14]
  PIN gpio_loopback_zero[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.490 4766.350 2881.790 4768.630 ;
    END
  END gpio_loopback_zero[15]
  PIN gpio_loopback_zero[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.490 4766.350 2384.790 4768.630 ;
    END
  END gpio_loopback_zero[16]
  PIN gpio_loopback_zero[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.490 4766.350 2128.790 4768.630 ;
    END
  END gpio_loopback_zero[17]
  PIN gpio_loopback_zero[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.490 4766.350 1683.790 4768.630 ;
    END
  END gpio_loopback_zero[18]
  PIN gpio_loopback_zero[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.490 4766.350 1161.790 4768.630 ;
    END
  END gpio_loopback_zero[19]
  PIN gpio_loopback_zero[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 615.030 3168.630 615.340 ;
    END
  END gpio_loopback_zero[1]
  PIN gpio_loopback_zero[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.490 4766.350 905.790 4768.630 ;
    END
  END gpio_loopback_zero[20]
  PIN gpio_loopback_zero[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.490 4766.350 649.790 4768.630 ;
    END
  END gpio_loopback_zero[21]
  PIN gpio_loopback_zero[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.490 4766.350 393.790 4768.630 ;
    END
  END gpio_loopback_zero[22]
  PIN gpio_loopback_zero[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.490 4766.350 137.790 4768.630 ;
    END
  END gpio_loopback_zero[23]
  PIN gpio_loopback_zero[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4523.220 0.300 4523.520 ;
    END
  END gpio_loopback_zero[24]
  PIN gpio_loopback_zero[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3673.220 0.300 3673.520 ;
    END
  END gpio_loopback_zero[25]
  PIN gpio_loopback_zero[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3458.220 0.300 3458.520 ;
    END
  END gpio_loopback_zero[26]
  PIN gpio_loopback_zero[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3243.220 0.300 3243.520 ;
    END
  END gpio_loopback_zero[27]
  PIN gpio_loopback_zero[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3028.220 0.300 3028.520 ;
    END
  END gpio_loopback_zero[28]
  PIN gpio_loopback_zero[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2813.220 0.300 2813.520 ;
    END
  END gpio_loopback_zero[29]
  PIN gpio_loopback_zero[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 840.030 3168.630 840.340 ;
    END
  END gpio_loopback_zero[2]
  PIN gpio_loopback_zero[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2598.220 0.300 2598.520 ;
    END
  END gpio_loopback_zero[30]
  PIN gpio_loopback_zero[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2383.220 0.300 2383.520 ;
    END
  END gpio_loopback_zero[31]
  PIN gpio_loopback_zero[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1738.220 0.300 1738.520 ;
    END
  END gpio_loopback_zero[32]
  PIN gpio_loopback_zero[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1523.220 0.300 1523.520 ;
    END
  END gpio_loopback_zero[33]
  PIN gpio_loopback_zero[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1308.220 0.300 1308.520 ;
    END
  END gpio_loopback_zero[34]
  PIN gpio_loopback_zero[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1093.220 0.300 1093.520 ;
    END
  END gpio_loopback_zero[35]
  PIN gpio_loopback_zero[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 878.220 0.300 878.520 ;
    END
  END gpio_loopback_zero[36]
  PIN gpio_loopback_zero[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 663.220 0.300 663.520 ;
    END
  END gpio_loopback_zero[37]
  PIN gpio_loopback_zero[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.955 -2.000 819.215 0.280 ;
    END
  END gpio_loopback_zero[38]
  PIN gpio_loopback_zero[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.800 -2.000 1367.060 0.280 ;
    END
  END gpio_loopback_zero[39]
  PIN gpio_loopback_zero[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1065.030 3168.630 1065.340 ;
    END
  END gpio_loopback_zero[3]
  PIN gpio_loopback_zero[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.825 -2.000 1641.085 0.280 ;
    END
  END gpio_loopback_zero[40]
  PIN gpio_loopback_zero[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.890 -2.000 1915.150 0.280 ;
    END
  END gpio_loopback_zero[41]
  PIN gpio_loopback_zero[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.890 -2.000 2189.150 0.280 ;
    END
  END gpio_loopback_zero[42]
  PIN gpio_loopback_zero[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.175 -2.000 2463.435 0.280 ;
    END
  END gpio_loopback_zero[43]
  PIN gpio_loopback_zero[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1290.030 3168.630 1290.340 ;
    END
  END gpio_loopback_zero[4]
  PIN gpio_loopback_zero[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1515.030 3168.630 1515.340 ;
    END
  END gpio_loopback_zero[5]
  PIN gpio_loopback_zero[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1740.030 3168.630 1740.340 ;
    END
  END gpio_loopback_zero[6]
  PIN gpio_loopback_zero[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2625.030 3168.630 2625.340 ;
    END
  END gpio_loopback_zero[7]
  PIN gpio_loopback_zero[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2850.030 3168.630 2850.340 ;
    END
  END gpio_loopback_zero[8]
  PIN gpio_loopback_zero[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3075.030 3168.630 3075.340 ;
    END
  END gpio_loopback_zero[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 364.760 3168.630 365.110 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3280.760 3168.630 3281.110 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3505.760 3168.630 3506.110 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3730.760 3168.630 3731.110 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4176.760 3168.630 4177.110 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4622.760 3168.630 4623.110 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2923.560 4766.350 2923.840 4768.630 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.560 4766.350 2414.840 4768.630 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.560 4766.350 2157.840 4768.630 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.560 4766.350 1712.840 4768.630 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.560 4766.350 1203.840 4768.630 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 590.760 3168.630 591.110 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.560 4766.350 945.840 4768.630 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.560 4766.350 688.840 4768.630 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.560 4766.350 431.840 4768.630 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.560 4766.350 174.840 4768.630 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4564.520 0.300 4564.870 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3715.520 0.300 3715.870 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3499.520 0.300 3499.870 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3283.520 0.300 3283.870 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3067.520 0.300 3067.870 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2851.520 0.300 2851.870 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 815.760 3168.630 816.110 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2635.520 0.300 2635.870 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2419.520 0.300 2419.870 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1781.520 0.300 1781.870 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1565.520 0.300 1565.870 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1349.520 0.300 1349.870 ;
    END
  END gpio_oeb[34]
  PIN gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1133.520 0.300 1133.870 ;
    END
  END gpio_oeb[35]
  PIN gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 917.520 0.300 917.870 ;
    END
  END gpio_oeb[36]
  PIN gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 701.520 0.300 701.870 ;
    END
  END gpio_oeb[37]
  PIN gpio_oeb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.790 -2.000 797.070 0.280 ;
    END
  END gpio_oeb[38]
  PIN gpio_oeb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.790 -2.000 1340.070 0.280 ;
    END
  END gpio_oeb[39]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1041.760 3168.630 1042.110 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.790 -2.000 1614.070 0.280 ;
    END
  END gpio_oeb[40]
  PIN gpio_oeb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -2.000 1888.070 0.280 ;
    END
  END gpio_oeb[41]
  PIN gpio_oeb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.790 -2.000 2162.070 0.280 ;
    END
  END gpio_oeb[42]
  PIN gpio_oeb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2435.790 -2.000 2436.070 0.280 ;
    END
  END gpio_oeb[43]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1266.760 3168.630 1267.110 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1491.760 3168.630 1492.110 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1717.760 3168.630 1718.110 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2603.760 3168.630 2604.110 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2829.760 3168.630 2830.110 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3054.760 3168.630 3055.110 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 349.120 3168.630 349.470 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3265.120 3168.630 3265.470 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3490.120 3168.630 3490.470 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3715.120 3168.630 3715.470 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4161.120 3168.630 4161.470 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4607.120 3168.630 4607.470 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2939.200 4766.350 2939.480 4768.630 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2430.200 4766.350 2430.480 4768.630 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.200 4766.350 2173.480 4768.630 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.200 4766.350 1728.480 4768.630 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.200 4766.350 1219.480 4768.630 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 575.120 3168.630 575.470 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.200 4766.350 961.480 4768.630 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.200 4766.350 704.480 4768.630 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.200 4766.350 447.480 4768.630 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.200 4766.350 190.480 4768.630 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4580.160 0.300 4580.510 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3731.160 0.300 3731.510 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3515.160 0.300 3515.510 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3299.160 0.300 3299.510 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3083.160 0.300 3083.510 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2867.160 0.300 2867.510 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 800.120 3168.630 800.470 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2651.160 0.300 2651.510 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2435.160 0.300 2435.510 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1797.160 0.300 1797.510 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1581.160 0.300 1581.510 ;
    END
  END gpio_out[33]
  PIN gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1365.160 0.300 1365.510 ;
    END
  END gpio_out[34]
  PIN gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1149.160 0.300 1149.510 ;
    END
  END gpio_out[35]
  PIN gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 933.160 0.300 933.510 ;
    END
  END gpio_out[36]
  PIN gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 717.160 0.300 717.510 ;
    END
  END gpio_out[37]
  PIN gpio_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.150 -2.000 781.430 0.280 ;
    END
  END gpio_out[38]
  PIN gpio_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.150 -2.000 1324.430 0.280 ;
    END
  END gpio_out[39]
  PIN gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1026.120 3168.630 1026.470 ;
    END
  END gpio_out[3]
  PIN gpio_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.150 -2.000 1598.430 0.280 ;
    END
  END gpio_out[40]
  PIN gpio_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.150 -2.000 1872.430 0.280 ;
    END
  END gpio_out[41]
  PIN gpio_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.150 -2.000 2146.430 0.280 ;
    END
  END gpio_out[42]
  PIN gpio_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.150 -2.000 2420.430 0.280 ;
    END
  END gpio_out[43]
  PIN gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1251.120 3168.630 1251.470 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1476.120 3168.630 1476.470 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1702.120 3168.630 1702.470 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2588.120 3168.630 2588.470 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2814.120 3168.630 2814.470 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3039.120 3168.630 3039.470 ;
    END
  END gpio_out[9]
  PIN gpio_slow_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 303.120 3168.630 303.470 ;
    END
  END gpio_slow_sel[0]
  PIN gpio_slow_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3219.120 3168.630 3219.470 ;
    END
  END gpio_slow_sel[10]
  PIN gpio_slow_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3444.120 3168.630 3444.470 ;
    END
  END gpio_slow_sel[11]
  PIN gpio_slow_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3669.120 3168.630 3669.470 ;
    END
  END gpio_slow_sel[12]
  PIN gpio_slow_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4115.120 3168.630 4115.470 ;
    END
  END gpio_slow_sel[13]
  PIN gpio_slow_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4561.120 3168.630 4561.470 ;
    END
  END gpio_slow_sel[14]
  PIN gpio_slow_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2985.200 4766.350 2985.480 4768.630 ;
    END
  END gpio_slow_sel[15]
  PIN gpio_slow_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.200 4766.350 2476.480 4768.630 ;
    END
  END gpio_slow_sel[16]
  PIN gpio_slow_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.200 4766.350 2219.480 4768.630 ;
    END
  END gpio_slow_sel[17]
  PIN gpio_slow_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.200 4766.350 1774.480 4768.630 ;
    END
  END gpio_slow_sel[18]
  PIN gpio_slow_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.200 4766.350 1265.480 4768.630 ;
    END
  END gpio_slow_sel[19]
  PIN gpio_slow_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 529.120 3168.630 529.470 ;
    END
  END gpio_slow_sel[1]
  PIN gpio_slow_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.200 4766.350 1007.480 4768.630 ;
    END
  END gpio_slow_sel[20]
  PIN gpio_slow_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.200 4766.350 750.480 4768.630 ;
    END
  END gpio_slow_sel[21]
  PIN gpio_slow_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.200 4766.350 493.480 4768.630 ;
    END
  END gpio_slow_sel[22]
  PIN gpio_slow_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.200 4766.350 236.480 4768.630 ;
    END
  END gpio_slow_sel[23]
  PIN gpio_slow_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4626.160 0.300 4626.510 ;
    END
  END gpio_slow_sel[24]
  PIN gpio_slow_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3777.160 0.300 3777.510 ;
    END
  END gpio_slow_sel[25]
  PIN gpio_slow_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3561.160 0.300 3561.510 ;
    END
  END gpio_slow_sel[26]
  PIN gpio_slow_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3345.160 0.300 3345.510 ;
    END
  END gpio_slow_sel[27]
  PIN gpio_slow_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3129.160 0.300 3129.510 ;
    END
  END gpio_slow_sel[28]
  PIN gpio_slow_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2913.160 0.300 2913.510 ;
    END
  END gpio_slow_sel[29]
  PIN gpio_slow_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 754.120 3168.630 754.470 ;
    END
  END gpio_slow_sel[2]
  PIN gpio_slow_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2697.160 0.300 2697.510 ;
    END
  END gpio_slow_sel[30]
  PIN gpio_slow_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2481.160 0.300 2481.510 ;
    END
  END gpio_slow_sel[31]
  PIN gpio_slow_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1843.160 0.300 1843.510 ;
    END
  END gpio_slow_sel[32]
  PIN gpio_slow_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1627.160 0.300 1627.510 ;
    END
  END gpio_slow_sel[33]
  PIN gpio_slow_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1411.160 0.300 1411.510 ;
    END
  END gpio_slow_sel[34]
  PIN gpio_slow_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1195.160 0.300 1195.510 ;
    END
  END gpio_slow_sel[35]
  PIN gpio_slow_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 979.160 0.300 979.510 ;
    END
  END gpio_slow_sel[36]
  PIN gpio_slow_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 763.160 0.300 763.510 ;
    END
  END gpio_slow_sel[37]
  PIN gpio_slow_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.150 -2.000 735.430 0.280 ;
    END
  END gpio_slow_sel[38]
  PIN gpio_slow_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.150 -2.000 1278.430 0.280 ;
    END
  END gpio_slow_sel[39]
  PIN gpio_slow_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 980.120 3168.630 980.470 ;
    END
  END gpio_slow_sel[3]
  PIN gpio_slow_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.150 -2.000 1552.430 0.280 ;
    END
  END gpio_slow_sel[40]
  PIN gpio_slow_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.150 -2.000 1826.430 0.280 ;
    END
  END gpio_slow_sel[41]
  PIN gpio_slow_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.150 -2.000 2100.430 0.280 ;
    END
  END gpio_slow_sel[42]
  PIN gpio_slow_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.150 -2.000 2374.430 0.280 ;
    END
  END gpio_slow_sel[43]
  PIN gpio_slow_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1205.120 3168.630 1205.470 ;
    END
  END gpio_slow_sel[4]
  PIN gpio_slow_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1430.120 3168.630 1430.470 ;
    END
  END gpio_slow_sel[5]
  PIN gpio_slow_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1656.120 3168.630 1656.470 ;
    END
  END gpio_slow_sel[6]
  PIN gpio_slow_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2542.120 3168.630 2542.470 ;
    END
  END gpio_slow_sel[7]
  PIN gpio_slow_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2768.120 3168.630 2768.470 ;
    END
  END gpio_slow_sel[8]
  PIN gpio_slow_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2993.120 3168.630 2993.470 ;
    END
  END gpio_slow_sel[9]
  PIN gpio_vtrip_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 358.320 3168.630 358.670 ;
    END
  END gpio_vtrip_sel[0]
  PIN gpio_vtrip_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3274.320 3168.630 3274.670 ;
    END
  END gpio_vtrip_sel[10]
  PIN gpio_vtrip_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3499.320 3168.630 3499.670 ;
    END
  END gpio_vtrip_sel[11]
  PIN gpio_vtrip_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3724.320 3168.630 3724.670 ;
    END
  END gpio_vtrip_sel[12]
  PIN gpio_vtrip_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4170.320 3168.630 4170.670 ;
    END
  END gpio_vtrip_sel[13]
  PIN gpio_vtrip_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4616.320 3168.630 4616.670 ;
    END
  END gpio_vtrip_sel[14]
  PIN gpio_vtrip_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2930.000 4766.350 2930.280 4768.630 ;
    END
  END gpio_vtrip_sel[15]
  PIN gpio_vtrip_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2421.000 4766.350 2421.280 4768.630 ;
    END
  END gpio_vtrip_sel[16]
  PIN gpio_vtrip_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.000 4766.350 2164.280 4768.630 ;
    END
  END gpio_vtrip_sel[17]
  PIN gpio_vtrip_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.000 4766.350 1719.280 4768.630 ;
    END
  END gpio_vtrip_sel[18]
  PIN gpio_vtrip_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.000 4766.350 1210.280 4768.630 ;
    END
  END gpio_vtrip_sel[19]
  PIN gpio_vtrip_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 584.320 3168.630 584.670 ;
    END
  END gpio_vtrip_sel[1]
  PIN gpio_vtrip_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.000 4766.350 952.280 4768.630 ;
    END
  END gpio_vtrip_sel[20]
  PIN gpio_vtrip_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.000 4766.350 695.280 4768.630 ;
    END
  END gpio_vtrip_sel[21]
  PIN gpio_vtrip_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.000 4766.350 438.280 4768.630 ;
    END
  END gpio_vtrip_sel[22]
  PIN gpio_vtrip_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.000 4766.350 181.280 4768.630 ;
    END
  END gpio_vtrip_sel[23]
  PIN gpio_vtrip_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 4570.960 0.300 4571.310 ;
    END
  END gpio_vtrip_sel[24]
  PIN gpio_vtrip_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3721.960 0.300 3722.310 ;
    END
  END gpio_vtrip_sel[25]
  PIN gpio_vtrip_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3505.960 0.300 3506.310 ;
    END
  END gpio_vtrip_sel[26]
  PIN gpio_vtrip_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3289.960 0.300 3290.310 ;
    END
  END gpio_vtrip_sel[27]
  PIN gpio_vtrip_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 3073.960 0.300 3074.310 ;
    END
  END gpio_vtrip_sel[28]
  PIN gpio_vtrip_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2857.960 0.300 2858.310 ;
    END
  END gpio_vtrip_sel[29]
  PIN gpio_vtrip_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 809.320 3168.630 809.670 ;
    END
  END gpio_vtrip_sel[2]
  PIN gpio_vtrip_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2641.960 0.300 2642.310 ;
    END
  END gpio_vtrip_sel[30]
  PIN gpio_vtrip_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2425.960 0.300 2426.310 ;
    END
  END gpio_vtrip_sel[31]
  PIN gpio_vtrip_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1787.960 0.300 1788.310 ;
    END
  END gpio_vtrip_sel[32]
  PIN gpio_vtrip_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1571.960 0.300 1572.310 ;
    END
  END gpio_vtrip_sel[33]
  PIN gpio_vtrip_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1355.960 0.300 1356.310 ;
    END
  END gpio_vtrip_sel[34]
  PIN gpio_vtrip_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1139.960 0.300 1140.310 ;
    END
  END gpio_vtrip_sel[35]
  PIN gpio_vtrip_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 923.960 0.300 924.310 ;
    END
  END gpio_vtrip_sel[36]
  PIN gpio_vtrip_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 707.960 0.300 708.310 ;
    END
  END gpio_vtrip_sel[37]
  PIN gpio_vtrip_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.350 -2.000 790.630 0.280 ;
    END
  END gpio_vtrip_sel[38]
  PIN gpio_vtrip_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.350 -2.000 1333.630 0.280 ;
    END
  END gpio_vtrip_sel[39]
  PIN gpio_vtrip_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1035.320 3168.630 1035.670 ;
    END
  END gpio_vtrip_sel[3]
  PIN gpio_vtrip_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.350 -2.000 1607.630 0.280 ;
    END
  END gpio_vtrip_sel[40]
  PIN gpio_vtrip_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.350 -2.000 1881.630 0.280 ;
    END
  END gpio_vtrip_sel[41]
  PIN gpio_vtrip_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.350 -2.000 2155.630 0.280 ;
    END
  END gpio_vtrip_sel[42]
  PIN gpio_vtrip_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.350 -2.000 2429.630 0.280 ;
    END
  END gpio_vtrip_sel[43]
  PIN gpio_vtrip_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1260.320 3168.630 1260.670 ;
    END
  END gpio_vtrip_sel[4]
  PIN gpio_vtrip_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1485.320 3168.630 1485.670 ;
    END
  END gpio_vtrip_sel[5]
  PIN gpio_vtrip_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1711.320 3168.630 1711.670 ;
    END
  END gpio_vtrip_sel[6]
  PIN gpio_vtrip_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2597.320 3168.630 2597.670 ;
    END
  END gpio_vtrip_sel[7]
  PIN gpio_vtrip_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2823.320 3168.630 2823.670 ;
    END
  END gpio_vtrip_sel[8]
  PIN gpio_vtrip_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3048.320 3168.630 3048.670 ;
    END
  END gpio_vtrip_sel[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3025.410 -2.000 3025.670 0.280 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3036.610 -2.000 3036.870 0.280 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3037.730 -2.000 3037.990 0.280 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3038.850 -2.000 3039.110 0.280 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3039.970 -2.000 3040.230 0.280 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3041.090 -2.000 3041.350 0.280 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3042.210 -2.000 3042.470 0.280 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3043.330 -2.000 3043.590 0.280 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3044.450 -2.000 3044.710 0.280 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3045.570 -2.000 3045.830 0.280 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3046.690 -2.000 3046.950 0.280 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3026.530 -2.000 3026.790 0.280 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3047.810 -2.000 3048.070 0.280 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3048.930 -2.000 3049.190 0.280 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3050.050 -2.000 3050.310 0.280 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3051.170 -2.000 3051.430 0.280 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3052.290 -2.000 3052.550 0.280 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3053.410 -2.000 3053.670 0.280 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3054.530 -2.000 3054.790 0.280 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3055.650 -2.000 3055.910 0.280 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3056.770 -2.000 3057.030 0.280 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3057.890 -2.000 3058.150 0.280 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3027.650 -2.000 3027.910 0.280 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3059.010 -2.000 3059.270 0.280 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3060.130 -2.000 3060.390 0.280 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3028.770 -2.000 3029.030 0.280 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3029.890 -2.000 3030.150 0.280 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3031.010 -2.000 3031.270 0.280 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3032.130 -2.000 3032.390 0.280 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3033.250 -2.000 3033.510 0.280 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3034.370 -2.000 3034.630 0.280 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3035.490 -2.000 3035.750 0.280 ;
    END
  END mask_rev[9]
  PIN por_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 266.860 0.300 267.210 ;
    END
  END por_l
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 265.735 0.300 266.085 ;
    END
  END porb_h
  PIN porb_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 267.975 0.300 268.325 ;
    END
  END porb_l
  PIN resetb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.880 -2.000 498.160 0.280 ;
    END
  END resetb_h
  PIN resetb_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.820 -2.000 551.100 0.280 ;
    END
  END resetb_l
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 129.810 0.300 153.810 ;
    END
  END vccd
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 180.070 0.300 204.020 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4327.610 3168.630 4351.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4377.810 3168.630 4401.810 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2114.050 3168.630 2137.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.020 24.800 44.020 4740.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 24.020 24.800 3142.620 44.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 24.020 4720.640 3142.620 4740.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 3122.620 24.800 3142.620 4740.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.250 2.400 61.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.250 2.400 101.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.250 2.400 141.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.250 2.400 181.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 215.250 2.400 221.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 255.250 2.400 261.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.250 2.400 301.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.250 2.400 341.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.250 2.400 381.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 415.250 2.400 421.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 455.250 2.400 461.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.250 2.400 501.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.250 2.400 541.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.250 2.400 581.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 615.250 2.400 621.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.250 2.400 661.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 695.250 2.400 701.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.250 2.400 741.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.250 2.400 781.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.250 2.400 821.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.250 2.400 861.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 895.250 2.400 901.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.250 2.400 941.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.250 2.400 981.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.250 2.400 1021.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.250 2.400 1061.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.250 2.400 1101.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.250 2.400 1141.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1175.250 2.400 1181.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.250 2.400 1221.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1255.250 2.400 1261.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.250 2.400 1301.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.250 2.400 1341.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.250 2.400 1381.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.250 2.400 1421.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1455.250 2.400 1461.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.250 2.400 1501.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.250 2.400 1541.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.250 2.400 1581.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1615.250 2.400 1621.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.250 2.400 1661.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1695.250 2.400 1701.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.250 2.400 1741.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.250 2.400 1781.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1815.250 2.400 1821.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1855.250 2.400 1861.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1895.250 2.400 1901.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.250 2.400 1941.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1975.250 2.400 1981.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2015.250 2.400 2021.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.250 2.400 2061.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2095.250 2.400 2101.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.250 2.400 2141.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.250 2.400 2181.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.250 2.400 2221.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.250 2.400 2261.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.250 2.400 2301.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2335.250 2.400 2341.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.250 2.400 2381.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2415.250 2.400 2421.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2455.250 2.400 2461.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2495.250 2.400 2501.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2535.250 2.400 2541.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2575.250 2.400 2581.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2615.250 2.400 2621.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.250 2.400 2661.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2695.250 2.400 2701.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.250 2.400 2741.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2775.250 2.400 2781.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2815.250 2.400 2821.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2855.250 2.400 2861.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2895.250 2.400 2901.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2935.250 2.400 2941.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2975.250 2.400 2981.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3015.250 2.400 3021.650 1472.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 3015.250 2213.445 3021.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3055.250 2.400 3061.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3095.250 2.400 3101.650 4763.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 60.430 3165.020 66.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 100.430 3165.020 106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 140.430 3165.020 146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 180.430 3165.020 186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 220.430 3165.020 226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 260.430 3165.020 266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 300.430 3165.020 306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 340.430 3165.020 346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 380.430 3165.020 386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 420.430 3165.020 426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 460.430 3165.020 466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 500.430 3165.020 506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 540.430 3165.020 546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 580.430 3165.020 586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 620.430 3165.020 626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 660.430 3165.020 666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 700.430 3165.020 706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 740.430 3165.020 746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 780.430 3165.020 786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 820.430 3165.020 826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 860.430 3165.020 866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 900.430 3165.020 906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 940.430 3165.020 946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 980.430 3165.020 986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1020.430 3165.020 1026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1060.430 3165.020 1066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1100.430 3165.020 1106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1140.430 3165.020 1146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1180.430 3165.020 1186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1220.430 3165.020 1226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1260.430 3165.020 1266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1300.430 3165.020 1306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1340.430 3165.020 1346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1380.430 3165.020 1386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1420.430 3165.020 1426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1460.430 3165.020 1466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1500.430 3165.020 1506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1540.430 3165.020 1546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1580.430 3165.020 1586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1620.430 3165.020 1626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1660.430 3165.020 1666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1700.430 3165.020 1706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1740.430 3165.020 1746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1780.430 3165.020 1786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1820.430 3165.020 1826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1860.430 3165.020 1866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1900.430 3165.020 1906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1940.430 3165.020 1946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1980.430 3165.020 1986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2020.430 3165.020 2026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2060.430 3165.020 2066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2100.430 3165.020 2106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2140.430 3165.020 2146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2180.430 3165.020 2186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2220.430 3165.020 2226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2260.430 3165.020 2266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2300.430 3165.020 2306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2340.430 3165.020 2346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2380.430 3165.020 2386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2420.430 3165.020 2426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2460.430 3165.020 2466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2500.430 3165.020 2506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2540.430 3165.020 2546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2580.430 3165.020 2586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2620.430 3165.020 2626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2660.430 3165.020 2666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2700.430 3165.020 2706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2740.430 3165.020 2746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2780.430 3165.020 2786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2820.430 3165.020 2826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2860.430 3165.020 2866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2900.430 3165.020 2906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2940.430 3165.020 2946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2980.430 3165.020 2986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3020.430 3165.020 3026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3060.430 3165.020 3066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3100.430 3165.020 3106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3140.430 3165.020 3146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3180.430 3165.020 3186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3220.430 3165.020 3226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3260.430 3165.020 3266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3300.430 3165.020 3306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3340.430 3165.020 3346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3380.430 3165.020 3386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3420.430 3165.020 3426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3460.430 3165.020 3466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3500.430 3165.020 3506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3540.430 3165.020 3546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3580.430 3165.020 3586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3620.430 3165.020 3626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3660.430 3165.020 3666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3700.430 3165.020 3706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3740.430 3165.020 3746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3780.430 3165.020 3786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3820.430 3165.020 3826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3860.430 3165.020 3866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3900.430 3165.020 3906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3940.430 3165.020 3946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3980.430 3165.020 3986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4020.430 3165.020 4026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4060.430 3165.020 4066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4100.430 3165.020 4106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4140.430 3165.020 4146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4180.430 3165.020 4186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4220.430 3165.020 4226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4260.430 3165.020 4266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4300.430 3165.020 4306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4340.430 3165.020 4346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4380.430 3165.020 4386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4420.430 3165.020 4426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4460.430 3165.020 4466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4500.430 3165.020 4506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4540.430 3165.020 4546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4580.430 3165.020 4586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4620.430 3165.020 4626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4660.430 3165.020 4666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4700.430 3165.020 4706.830 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 2019.310 0.300 2042.570 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 4349.820 0.300 4373.820 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 4400.070 0.300 4424.020 ;
    END
  END vccd2
  PIN vdda
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2904.030 -2.000 2927.930 0.300 ;
    END
  END vdda
  PIN vdda
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2953.920 -2.000 2977.820 0.300 ;
    END
  END vdda
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3882.030 3168.630 3905.930 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2309.020 3168.630 2332.920 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2358.920 3168.630 2382.820 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 3166.330 3931.920 3168.630 3955.820 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 2254.700 0.300 2278.600 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 2204.810 0.300 2228.710 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 390.700 0.300 414.600 ;
    END
  END vddio
  PIN vddio
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 4188.710 0.300 4212.610 ;
    END
  END vddio
  PIN vddio
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 340.810 0.300 364.710 ;
    END
  END vddio
  PIN vddio
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -2.000 4138.810 0.300 4162.710 ;
    END
  END vddio
  PIN vssa
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 233.920 -2.000 257.820 0.300 ;
    END
  END vssa
  PIN vssa
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 184.030 -2.000 207.930 0.300 ;
    END
  END vssa
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2717.710 4766.330 2741.610 4768.630 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1868.030 3168.630 1891.930 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2667.810 4766.330 2691.710 4768.630 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3166.330 1917.920 3168.630 1941.820 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -2.000 3977.710 0.300 4001.610 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -2.000 3927.810 0.300 3951.710 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 1045.820 -2.000 1069.820 0.300 ;
    END
  END vssd
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 996.420 -2.000 1019.570 0.300 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3166.330 4353.050 3168.630 4376.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2138.810 3168.630 2162.810 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3166.330 2088.610 3168.630 2112.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.620 2.400 21.620 4763.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2.400 3165.020 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4743.040 3165.020 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3145.020 2.400 3165.020 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.850 2.400 71.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.850 2.400 111.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.850 2.400 151.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.850 2.400 191.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.850 2.400 231.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.850 2.400 271.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.850 2.400 311.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.850 2.400 351.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.850 2.400 391.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.850 2.400 431.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.850 2.400 471.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.850 2.400 511.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.850 2.400 551.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.850 2.400 591.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.850 2.400 631.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.850 2.400 671.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.850 2.400 711.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.850 2.400 751.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.850 2.400 791.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.850 2.400 831.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.850 2.400 871.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.850 2.400 911.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 944.850 2.400 951.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 984.850 2.400 991.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.850 2.400 1031.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.850 2.400 1071.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.850 2.400 1111.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.850 2.400 1151.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.850 2.400 1191.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.850 2.400 1231.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.850 2.400 1271.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.850 2.400 1311.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.850 2.400 1351.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1384.850 2.400 1391.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1424.850 2.400 1431.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.850 2.400 1471.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.850 2.400 1511.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.850 2.400 1551.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.850 2.400 1591.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1624.850 2.400 1631.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.850 2.400 1671.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.850 2.400 1711.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.850 2.400 1751.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1784.850 2.400 1791.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1824.850 2.400 1831.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.850 2.400 1871.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.850 2.400 1911.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1944.850 2.400 1951.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.850 2.400 1991.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.850 2.400 2031.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.850 2.400 2071.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.850 2.400 2111.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.850 2.400 2151.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.850 2.400 2191.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.850 2.400 2231.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.850 2.400 2271.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.850 2.400 2311.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.850 2.400 2351.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2384.850 2.400 2391.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.850 2.400 2431.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.850 2.400 2471.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.850 2.400 2511.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2544.850 2.400 2551.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.850 2.400 2591.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.850 2.400 2631.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.850 2.400 2671.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.850 2.400 2711.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2744.850 2.400 2751.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2784.850 2.400 2791.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2824.850 2.400 2831.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2864.850 2.400 2871.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2904.850 2.400 2911.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2944.850 2.400 2951.250 234.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2944.850 3732.980 2951.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2984.850 2.400 2991.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3024.850 2.400 3031.250 234.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 3024.850 3732.980 3031.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3064.850 2.400 3071.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3104.850 2.400 3111.250 4763.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 70.030 3165.020 76.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 110.030 3165.020 116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 150.030 3165.020 156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 190.030 3165.020 196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 230.030 3165.020 236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 270.030 3165.020 276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 310.030 3165.020 316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 350.030 3165.020 356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 390.030 3165.020 396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 430.030 3165.020 436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 470.030 3165.020 476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 510.030 3165.020 516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 550.030 3165.020 556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 590.030 3165.020 596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 630.030 3165.020 636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 670.030 3165.020 676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 710.030 3165.020 716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 750.030 3165.020 756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 790.030 3165.020 796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 830.030 3165.020 836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 870.030 3165.020 876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 910.030 3165.020 916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 950.030 3165.020 956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 990.030 3165.020 996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1030.030 3165.020 1036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1070.030 3165.020 1076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1110.030 3165.020 1116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1150.030 3165.020 1156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1190.030 3165.020 1196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1230.030 3165.020 1236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1270.030 3165.020 1276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1310.030 3165.020 1316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1350.030 3165.020 1356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1390.030 3165.020 1396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1430.030 3165.020 1436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1470.030 3165.020 1476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1510.030 3165.020 1516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1550.030 3165.020 1556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1590.030 3165.020 1596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1630.030 3165.020 1636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1670.030 3165.020 1676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1710.030 3165.020 1716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1750.030 3165.020 1756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1790.030 3165.020 1796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1830.030 3165.020 1836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1870.030 3165.020 1876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1910.030 3165.020 1916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1950.030 3165.020 1956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1990.030 3165.020 1996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2030.030 3165.020 2036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2070.030 3165.020 2076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2110.030 3165.020 2116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2150.030 3165.020 2156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2190.030 3165.020 2196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2230.030 3165.020 2236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2270.030 3165.020 2276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2310.030 3165.020 2316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2350.030 3165.020 2356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2390.030 3165.020 2396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2430.030 3165.020 2436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2470.030 3165.020 2476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2510.030 3165.020 2516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2550.030 3165.020 2556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2590.030 3165.020 2596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2630.030 3165.020 2636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2670.030 3165.020 2676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2710.030 3165.020 2716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2750.030 3165.020 2756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2790.030 3165.020 2796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2830.030 3165.020 2836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2870.030 3165.020 2876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2910.030 3165.020 2916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2950.030 3165.020 2956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2990.030 3165.020 2996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3030.030 3165.020 3036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3070.030 3165.020 3076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3110.030 3165.020 3116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3150.030 3165.020 3156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3190.030 3165.020 3196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3230.030 3165.020 3236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3270.030 3165.020 3276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3310.030 3165.020 3316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3350.030 3165.020 3356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3390.030 3165.020 3396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3430.030 3165.020 3436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3470.030 3165.020 3476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3510.030 3165.020 3516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3550.030 3165.020 3556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3590.030 3165.020 3596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3630.030 3165.020 3636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3670.030 3165.020 3676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3710.030 3165.020 3716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3750.030 3165.020 3756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3790.030 3165.020 3796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3830.030 3165.020 3836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3870.030 3165.020 3876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3910.030 3165.020 3916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3950.030 3165.020 3956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3990.030 3165.020 3996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4030.030 3165.020 4036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4070.030 3165.020 4076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4110.030 3165.020 4116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4150.030 3165.020 4156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4190.030 3165.020 4196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4230.030 3165.020 4236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4270.030 3165.020 4276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4310.030 3165.020 4316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4350.030 3165.020 4356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4390.030 3165.020 4396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4430.030 3165.020 4436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4470.030 3165.020 4476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4510.030 3165.020 4516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4550.030 3165.020 4556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4590.030 3165.020 4596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4630.030 3165.020 4636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4670.030 3165.020 4676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4710.030 3165.020 4716.430 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -2.000 1993.810 0.300 2017.810 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -2.000 2044.070 0.300 2068.020 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -2.000 4375.270 0.300 4398.580 ;
    END
  END vssd2
  PIN vssio
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2635.030 -2.000 2658.930 0.300 ;
    END
  END vssio
  PIN vssio
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 1506.710 4766.330 1530.610 4768.630 ;
    END
  END vssio
  PIN vssio
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2684.920 -2.000 2708.820 0.300 ;
    END
  END vssio
  PIN vssio
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 1456.810 4766.330 1480.710 4768.630 ;
    END
  END vssio
  OBS
      LAYER li1 ;
        RECT 2855.880 245.795 3044.480 3722.125 ;
      LAYER met1 ;
        RECT 198.790 0.040 3045.330 4766.420 ;
      LAYER met2 ;
        RECT 0.090 4766.070 137.210 4766.530 ;
        RECT 138.070 4766.070 147.210 4766.530 ;
        RECT 148.070 4766.070 171.520 4766.530 ;
        RECT 172.360 4766.070 174.280 4766.530 ;
        RECT 175.120 4766.070 177.500 4766.530 ;
        RECT 178.340 4766.070 180.720 4766.530 ;
        RECT 181.560 4766.070 189.920 4766.530 ;
        RECT 190.760 4766.070 192.680 4766.530 ;
        RECT 193.520 4766.070 195.900 4766.530 ;
        RECT 196.740 4766.070 199.120 4766.530 ;
        RECT 199.960 4766.070 211.540 4766.530 ;
        RECT 212.380 4766.070 214.300 4766.530 ;
        RECT 215.140 4766.070 217.520 4766.530 ;
        RECT 218.360 4766.070 220.740 4766.530 ;
        RECT 221.580 4766.070 223.105 4766.530 ;
        RECT 224.735 4766.070 226.720 4766.530 ;
        RECT 227.560 4766.070 232.520 4766.530 ;
        RECT 233.720 4766.070 235.920 4766.530 ;
        RECT 236.760 4766.070 245.120 4766.530 ;
        RECT 245.960 4766.070 393.210 4766.530 ;
        RECT 394.070 4766.070 403.210 4766.530 ;
        RECT 404.070 4766.070 428.520 4766.530 ;
        RECT 429.360 4766.070 431.280 4766.530 ;
        RECT 432.120 4766.070 434.500 4766.530 ;
        RECT 435.340 4766.070 437.720 4766.530 ;
        RECT 438.560 4766.070 446.920 4766.530 ;
        RECT 447.760 4766.070 449.680 4766.530 ;
        RECT 450.520 4766.070 452.900 4766.530 ;
        RECT 453.740 4766.070 456.120 4766.530 ;
        RECT 456.960 4766.070 468.540 4766.530 ;
        RECT 469.380 4766.070 471.300 4766.530 ;
        RECT 472.140 4766.070 474.520 4766.530 ;
        RECT 475.360 4766.070 477.740 4766.530 ;
        RECT 478.580 4766.070 480.105 4766.530 ;
        RECT 481.735 4766.070 483.720 4766.530 ;
        RECT 484.560 4766.070 489.520 4766.530 ;
        RECT 490.720 4766.070 492.920 4766.530 ;
        RECT 493.760 4766.070 502.120 4766.530 ;
        RECT 502.960 4766.070 649.210 4766.530 ;
        RECT 650.070 4766.070 659.210 4766.530 ;
        RECT 660.070 4766.070 685.520 4766.530 ;
        RECT 686.360 4766.070 688.280 4766.530 ;
        RECT 689.120 4766.070 691.500 4766.530 ;
        RECT 692.340 4766.070 694.720 4766.530 ;
        RECT 695.560 4766.070 703.920 4766.530 ;
        RECT 704.760 4766.070 706.680 4766.530 ;
        RECT 707.520 4766.070 709.900 4766.530 ;
        RECT 710.740 4766.070 713.120 4766.530 ;
        RECT 713.960 4766.070 725.540 4766.530 ;
        RECT 726.380 4766.070 728.300 4766.530 ;
        RECT 729.140 4766.070 731.520 4766.530 ;
        RECT 732.360 4766.070 734.740 4766.530 ;
        RECT 735.580 4766.070 737.105 4766.530 ;
        RECT 738.735 4766.070 740.720 4766.530 ;
        RECT 741.560 4766.070 746.520 4766.530 ;
        RECT 747.720 4766.070 749.920 4766.530 ;
        RECT 750.760 4766.070 759.120 4766.530 ;
        RECT 759.960 4766.070 905.210 4766.530 ;
        RECT 906.070 4766.070 915.210 4766.530 ;
        RECT 916.070 4766.070 942.520 4766.530 ;
        RECT 943.360 4766.070 945.280 4766.530 ;
        RECT 946.120 4766.070 948.500 4766.530 ;
        RECT 949.340 4766.070 951.720 4766.530 ;
        RECT 952.560 4766.070 960.920 4766.530 ;
        RECT 961.760 4766.070 963.680 4766.530 ;
        RECT 964.520 4766.070 966.900 4766.530 ;
        RECT 967.740 4766.070 970.120 4766.530 ;
        RECT 970.960 4766.070 982.540 4766.530 ;
        RECT 983.380 4766.070 985.300 4766.530 ;
        RECT 986.140 4766.070 988.520 4766.530 ;
        RECT 989.360 4766.070 991.740 4766.530 ;
        RECT 992.580 4766.070 994.105 4766.530 ;
        RECT 995.735 4766.070 997.720 4766.530 ;
        RECT 998.560 4766.070 1003.520 4766.530 ;
        RECT 1004.720 4766.070 1006.920 4766.530 ;
        RECT 1007.760 4766.070 1016.120 4766.530 ;
        RECT 1016.960 4766.070 1161.210 4766.530 ;
        RECT 1162.070 4766.070 1171.210 4766.530 ;
        RECT 1172.070 4766.070 1200.520 4766.530 ;
        RECT 1201.360 4766.070 1203.280 4766.530 ;
        RECT 1204.120 4766.070 1206.500 4766.530 ;
        RECT 1207.340 4766.070 1209.720 4766.530 ;
        RECT 1210.560 4766.070 1218.920 4766.530 ;
        RECT 1219.760 4766.070 1221.680 4766.530 ;
        RECT 1222.520 4766.070 1224.900 4766.530 ;
        RECT 1225.740 4766.070 1228.120 4766.530 ;
        RECT 1228.960 4766.070 1240.540 4766.530 ;
        RECT 1241.380 4766.070 1243.300 4766.530 ;
        RECT 1244.140 4766.070 1246.520 4766.530 ;
        RECT 1247.360 4766.070 1249.740 4766.530 ;
        RECT 1250.580 4766.070 1252.105 4766.530 ;
        RECT 1253.735 4766.070 1255.720 4766.530 ;
        RECT 1256.560 4766.070 1261.520 4766.530 ;
        RECT 1262.720 4766.070 1264.920 4766.530 ;
        RECT 1265.760 4766.070 1274.120 4766.530 ;
        RECT 1274.960 4766.070 1683.210 4766.530 ;
        RECT 1684.070 4766.070 1693.210 4766.530 ;
        RECT 1694.070 4766.070 1709.520 4766.530 ;
        RECT 1710.360 4766.070 1712.280 4766.530 ;
        RECT 1713.120 4766.070 1715.500 4766.530 ;
        RECT 1716.340 4766.070 1718.720 4766.530 ;
        RECT 1719.560 4766.070 1727.920 4766.530 ;
        RECT 1728.760 4766.070 1730.680 4766.530 ;
        RECT 1731.520 4766.070 1733.900 4766.530 ;
        RECT 1734.740 4766.070 1737.120 4766.530 ;
        RECT 1737.960 4766.070 1749.540 4766.530 ;
        RECT 1750.380 4766.070 1752.300 4766.530 ;
        RECT 1753.140 4766.070 1755.520 4766.530 ;
        RECT 1756.360 4766.070 1758.740 4766.530 ;
        RECT 1759.580 4766.070 1761.105 4766.530 ;
        RECT 1762.735 4766.070 1764.720 4766.530 ;
        RECT 1765.560 4766.070 1770.520 4766.530 ;
        RECT 1771.720 4766.070 1773.920 4766.530 ;
        RECT 1774.760 4766.070 1783.120 4766.530 ;
        RECT 1783.960 4766.070 2128.210 4766.530 ;
        RECT 2129.070 4766.070 2138.210 4766.530 ;
        RECT 2139.070 4766.070 2154.520 4766.530 ;
        RECT 2155.360 4766.070 2157.280 4766.530 ;
        RECT 2158.120 4766.070 2160.500 4766.530 ;
        RECT 2161.340 4766.070 2163.720 4766.530 ;
        RECT 2164.560 4766.070 2172.920 4766.530 ;
        RECT 2173.760 4766.070 2175.680 4766.530 ;
        RECT 2176.520 4766.070 2178.900 4766.530 ;
        RECT 2179.740 4766.070 2182.120 4766.530 ;
        RECT 2182.960 4766.070 2194.540 4766.530 ;
        RECT 2195.380 4766.070 2197.300 4766.530 ;
        RECT 2198.140 4766.070 2200.520 4766.530 ;
        RECT 2201.360 4766.070 2203.740 4766.530 ;
        RECT 2204.580 4766.070 2206.105 4766.530 ;
        RECT 2207.735 4766.070 2209.720 4766.530 ;
        RECT 2210.560 4766.070 2215.520 4766.530 ;
        RECT 2216.720 4766.070 2218.920 4766.530 ;
        RECT 2219.760 4766.070 2228.120 4766.530 ;
        RECT 2228.960 4766.070 2384.210 4766.530 ;
        RECT 2385.070 4766.070 2394.210 4766.530 ;
        RECT 2395.070 4766.070 2411.520 4766.530 ;
        RECT 2412.360 4766.070 2414.280 4766.530 ;
        RECT 2415.120 4766.070 2417.500 4766.530 ;
        RECT 2418.340 4766.070 2420.720 4766.530 ;
        RECT 2421.560 4766.070 2429.920 4766.530 ;
        RECT 2430.760 4766.070 2432.680 4766.530 ;
        RECT 2433.520 4766.070 2435.900 4766.530 ;
        RECT 2436.740 4766.070 2439.120 4766.530 ;
        RECT 2439.960 4766.070 2451.540 4766.530 ;
        RECT 2452.380 4766.070 2454.300 4766.530 ;
        RECT 2455.140 4766.070 2457.520 4766.530 ;
        RECT 2458.360 4766.070 2460.740 4766.530 ;
        RECT 2461.580 4766.070 2463.105 4766.530 ;
        RECT 2464.735 4766.070 2466.720 4766.530 ;
        RECT 2467.560 4766.070 2472.520 4766.530 ;
        RECT 2473.720 4766.070 2475.920 4766.530 ;
        RECT 2476.760 4766.070 2485.120 4766.530 ;
        RECT 2485.960 4766.070 2881.210 4766.530 ;
        RECT 2882.070 4766.070 2891.210 4766.530 ;
        RECT 2892.070 4766.070 2920.520 4766.530 ;
        RECT 2921.360 4766.070 2923.280 4766.530 ;
        RECT 2924.120 4766.070 2926.500 4766.530 ;
        RECT 2927.340 4766.070 2929.720 4766.530 ;
        RECT 2930.560 4766.070 2938.920 4766.530 ;
        RECT 2939.760 4766.070 2941.680 4766.530 ;
        RECT 2942.520 4766.070 2944.900 4766.530 ;
        RECT 2945.740 4766.070 2948.120 4766.530 ;
        RECT 2948.960 4766.070 2960.540 4766.530 ;
        RECT 2961.380 4766.070 2963.300 4766.530 ;
        RECT 2964.140 4766.070 2966.520 4766.530 ;
        RECT 2967.360 4766.070 2969.740 4766.530 ;
        RECT 2970.580 4766.070 2972.105 4766.530 ;
        RECT 2973.735 4766.070 2975.720 4766.530 ;
        RECT 2976.560 4766.070 2981.520 4766.530 ;
        RECT 2982.720 4766.070 2984.920 4766.530 ;
        RECT 2985.760 4766.070 2994.120 4766.530 ;
        RECT 2994.960 4766.070 3166.550 4766.530 ;
        RECT 0.090 0.560 3166.550 4766.070 ;
        RECT 0.090 0.010 497.600 0.560 ;
        RECT 498.440 0.010 550.540 0.560 ;
        RECT 551.380 0.010 725.670 0.560 ;
        RECT 726.510 0.010 734.870 0.560 ;
        RECT 735.710 0.010 737.910 0.560 ;
        RECT 739.110 0.010 744.070 0.560 ;
        RECT 744.910 0.010 746.895 0.560 ;
        RECT 748.525 0.010 750.050 0.560 ;
        RECT 750.890 0.010 753.270 0.560 ;
        RECT 754.110 0.010 756.490 0.560 ;
        RECT 757.330 0.010 759.250 0.560 ;
        RECT 760.090 0.010 771.670 0.560 ;
        RECT 772.510 0.010 774.890 0.560 ;
        RECT 775.730 0.010 778.110 0.560 ;
        RECT 778.950 0.010 780.870 0.560 ;
        RECT 781.710 0.010 790.070 0.560 ;
        RECT 790.910 0.010 793.290 0.560 ;
        RECT 794.130 0.010 796.510 0.560 ;
        RECT 797.350 0.010 799.270 0.560 ;
        RECT 800.110 0.010 802.620 0.560 ;
        RECT 803.440 0.010 818.675 0.560 ;
        RECT 819.495 0.010 1268.670 0.560 ;
        RECT 1269.510 0.010 1277.870 0.560 ;
        RECT 1278.710 0.010 1280.910 0.560 ;
        RECT 1282.110 0.010 1287.070 0.560 ;
        RECT 1287.910 0.010 1289.895 0.560 ;
        RECT 1291.525 0.010 1293.050 0.560 ;
        RECT 1293.890 0.010 1296.270 0.560 ;
        RECT 1297.110 0.010 1299.490 0.560 ;
        RECT 1300.330 0.010 1302.250 0.560 ;
        RECT 1303.090 0.010 1314.670 0.560 ;
        RECT 1315.510 0.010 1317.890 0.560 ;
        RECT 1318.730 0.010 1321.110 0.560 ;
        RECT 1321.950 0.010 1323.870 0.560 ;
        RECT 1324.710 0.010 1333.070 0.560 ;
        RECT 1333.910 0.010 1336.290 0.560 ;
        RECT 1337.130 0.010 1339.510 0.560 ;
        RECT 1340.350 0.010 1342.270 0.560 ;
        RECT 1343.110 0.010 1345.620 0.560 ;
        RECT 1346.440 0.010 1366.520 0.560 ;
        RECT 1367.340 0.010 1542.670 0.560 ;
        RECT 1543.510 0.010 1551.870 0.560 ;
        RECT 1552.710 0.010 1554.910 0.560 ;
        RECT 1556.110 0.010 1561.070 0.560 ;
        RECT 1561.910 0.010 1563.895 0.560 ;
        RECT 1565.525 0.010 1567.050 0.560 ;
        RECT 1567.890 0.010 1570.270 0.560 ;
        RECT 1571.110 0.010 1573.490 0.560 ;
        RECT 1574.330 0.010 1576.250 0.560 ;
        RECT 1577.090 0.010 1588.670 0.560 ;
        RECT 1589.510 0.010 1591.890 0.560 ;
        RECT 1592.730 0.010 1595.110 0.560 ;
        RECT 1595.950 0.010 1597.870 0.560 ;
        RECT 1598.710 0.010 1607.070 0.560 ;
        RECT 1607.910 0.010 1610.290 0.560 ;
        RECT 1611.130 0.010 1613.510 0.560 ;
        RECT 1614.350 0.010 1616.270 0.560 ;
        RECT 1617.110 0.010 1619.620 0.560 ;
        RECT 1620.440 0.010 1640.545 0.560 ;
        RECT 1641.365 0.010 1816.670 0.560 ;
        RECT 1817.510 0.010 1825.870 0.560 ;
        RECT 1826.710 0.010 1828.910 0.560 ;
        RECT 1830.110 0.010 1835.070 0.560 ;
        RECT 1835.910 0.010 1837.895 0.560 ;
        RECT 1839.525 0.010 1841.050 0.560 ;
        RECT 1841.890 0.010 1844.270 0.560 ;
        RECT 1845.110 0.010 1847.490 0.560 ;
        RECT 1848.330 0.010 1850.250 0.560 ;
        RECT 1851.090 0.010 1862.670 0.560 ;
        RECT 1863.510 0.010 1865.890 0.560 ;
        RECT 1866.730 0.010 1869.110 0.560 ;
        RECT 1869.950 0.010 1871.870 0.560 ;
        RECT 1872.710 0.010 1881.070 0.560 ;
        RECT 1881.910 0.010 1884.290 0.560 ;
        RECT 1885.130 0.010 1887.510 0.560 ;
        RECT 1888.350 0.010 1890.270 0.560 ;
        RECT 1891.110 0.010 1893.620 0.560 ;
        RECT 1894.440 0.010 1914.610 0.560 ;
        RECT 1915.430 0.010 2090.670 0.560 ;
        RECT 2091.510 0.010 2099.870 0.560 ;
        RECT 2100.710 0.010 2102.910 0.560 ;
        RECT 2104.110 0.010 2109.070 0.560 ;
        RECT 2109.910 0.010 2111.895 0.560 ;
        RECT 2113.525 0.010 2115.050 0.560 ;
        RECT 2115.890 0.010 2118.270 0.560 ;
        RECT 2119.110 0.010 2121.490 0.560 ;
        RECT 2122.330 0.010 2124.250 0.560 ;
        RECT 2125.090 0.010 2136.670 0.560 ;
        RECT 2137.510 0.010 2139.890 0.560 ;
        RECT 2140.730 0.010 2143.110 0.560 ;
        RECT 2143.950 0.010 2145.870 0.560 ;
        RECT 2146.710 0.010 2155.070 0.560 ;
        RECT 2155.910 0.010 2158.290 0.560 ;
        RECT 2159.130 0.010 2161.510 0.560 ;
        RECT 2162.350 0.010 2164.270 0.560 ;
        RECT 2165.110 0.010 2167.620 0.560 ;
        RECT 2168.440 0.010 2188.610 0.560 ;
        RECT 2189.430 0.010 2364.670 0.560 ;
        RECT 2365.510 0.010 2373.870 0.560 ;
        RECT 2374.710 0.010 2376.910 0.560 ;
        RECT 2378.110 0.010 2383.070 0.560 ;
        RECT 2383.910 0.010 2385.895 0.560 ;
        RECT 2387.525 0.010 2389.050 0.560 ;
        RECT 2389.890 0.010 2392.270 0.560 ;
        RECT 2393.110 0.010 2395.490 0.560 ;
        RECT 2396.330 0.010 2398.250 0.560 ;
        RECT 2399.090 0.010 2410.670 0.560 ;
        RECT 2411.510 0.010 2413.890 0.560 ;
        RECT 2414.730 0.010 2417.110 0.560 ;
        RECT 2417.950 0.010 2419.870 0.560 ;
        RECT 2420.710 0.010 2429.070 0.560 ;
        RECT 2429.910 0.010 2432.290 0.560 ;
        RECT 2433.130 0.010 2435.510 0.560 ;
        RECT 2436.350 0.010 2438.270 0.560 ;
        RECT 2439.110 0.010 2441.620 0.560 ;
        RECT 2442.440 0.010 2462.895 0.560 ;
        RECT 2463.715 0.010 3025.130 0.560 ;
        RECT 3025.950 0.010 3026.250 0.560 ;
        RECT 3027.070 0.010 3027.370 0.560 ;
        RECT 3028.190 0.010 3028.490 0.560 ;
        RECT 3029.310 0.010 3029.610 0.560 ;
        RECT 3030.430 0.010 3030.730 0.560 ;
        RECT 3031.550 0.010 3031.850 0.560 ;
        RECT 3032.670 0.010 3032.970 0.560 ;
        RECT 3033.790 0.010 3034.090 0.560 ;
        RECT 3034.910 0.010 3035.210 0.560 ;
        RECT 3036.030 0.010 3036.330 0.560 ;
        RECT 3037.150 0.010 3037.450 0.560 ;
        RECT 3038.270 0.010 3038.570 0.560 ;
        RECT 3039.390 0.010 3039.690 0.560 ;
        RECT 3040.510 0.010 3040.810 0.560 ;
        RECT 3041.630 0.010 3041.930 0.560 ;
        RECT 3042.750 0.010 3043.050 0.560 ;
        RECT 3043.870 0.010 3044.170 0.560 ;
        RECT 3044.990 0.010 3045.290 0.560 ;
        RECT 3046.110 0.010 3046.410 0.560 ;
        RECT 3047.230 0.010 3047.530 0.560 ;
        RECT 3048.350 0.010 3048.650 0.560 ;
        RECT 3049.470 0.010 3049.770 0.560 ;
        RECT 3050.590 0.010 3050.890 0.560 ;
        RECT 3051.710 0.010 3052.010 0.560 ;
        RECT 3052.830 0.010 3053.130 0.560 ;
        RECT 3053.950 0.010 3054.250 0.560 ;
        RECT 3055.070 0.010 3055.370 0.560 ;
        RECT 3056.190 0.010 3056.490 0.560 ;
        RECT 3057.310 0.010 3057.610 0.560 ;
        RECT 3058.430 0.010 3058.730 0.560 ;
        RECT 3059.550 0.010 3059.850 0.560 ;
        RECT 3060.670 0.010 3166.550 0.560 ;
      LAYER met3 ;
        RECT 0.000 4645.740 3166.630 4746.905 ;
        RECT 0.000 4644.630 3165.930 4645.740 ;
        RECT 0.000 4636.110 3166.630 4644.630 ;
        RECT 0.700 4635.740 3166.630 4636.110 ;
        RECT 0.700 4634.960 3165.930 4635.740 ;
        RECT 0.000 4634.630 3165.930 4634.960 ;
        RECT 0.000 4626.910 3166.630 4634.630 ;
        RECT 0.700 4626.270 3166.630 4626.910 ;
        RECT 0.700 4625.760 3165.930 4626.270 ;
        RECT 0.000 4625.120 3165.930 4625.760 ;
        RECT 0.000 4623.840 3166.630 4625.120 ;
        RECT 0.700 4623.510 3166.630 4623.840 ;
        RECT 0.700 4622.400 3165.930 4623.510 ;
        RECT 0.000 4622.360 3165.930 4622.400 ;
        RECT 0.000 4620.290 3166.630 4622.360 ;
        RECT 0.000 4619.140 3165.930 4620.290 ;
        RECT 0.000 4617.710 3166.630 4619.140 ;
        RECT 0.700 4617.070 3166.630 4617.710 ;
        RECT 0.700 4616.560 3165.930 4617.070 ;
        RECT 0.000 4615.920 3165.930 4616.560 ;
        RECT 0.000 4614.855 3166.630 4615.920 ;
        RECT 0.700 4612.985 3166.630 4614.855 ;
        RECT 0.000 4611.730 3166.630 4612.985 ;
        RECT 0.700 4610.580 3166.630 4611.730 ;
        RECT 0.000 4608.510 3166.630 4610.580 ;
        RECT 0.700 4607.870 3166.630 4608.510 ;
        RECT 0.700 4607.360 3165.930 4607.870 ;
        RECT 0.000 4606.720 3165.930 4607.360 ;
        RECT 0.000 4605.290 3166.630 4606.720 ;
        RECT 0.700 4605.110 3166.630 4605.290 ;
        RECT 0.700 4604.140 3165.930 4605.110 ;
        RECT 0.000 4603.960 3165.930 4604.140 ;
        RECT 0.000 4602.530 3166.630 4603.960 ;
        RECT 0.700 4601.890 3166.630 4602.530 ;
        RECT 0.700 4601.380 3165.930 4601.890 ;
        RECT 0.000 4600.740 3165.930 4601.380 ;
        RECT 0.000 4598.670 3166.630 4600.740 ;
        RECT 0.000 4597.520 3165.930 4598.670 ;
        RECT 0.000 4590.110 3166.630 4597.520 ;
        RECT 0.700 4588.960 3166.630 4590.110 ;
        RECT 0.000 4586.890 3166.630 4588.960 ;
        RECT 0.700 4586.250 3166.630 4586.890 ;
        RECT 0.700 4585.740 3165.930 4586.250 ;
        RECT 0.000 4585.100 3165.930 4585.740 ;
        RECT 0.000 4583.670 3166.630 4585.100 ;
        RECT 0.700 4583.490 3166.630 4583.670 ;
        RECT 0.700 4582.520 3165.930 4583.490 ;
        RECT 0.000 4582.340 3165.930 4582.520 ;
        RECT 0.000 4580.910 3166.630 4582.340 ;
        RECT 0.700 4580.270 3166.630 4580.910 ;
        RECT 0.700 4579.760 3165.930 4580.270 ;
        RECT 0.000 4579.120 3165.930 4579.760 ;
        RECT 0.000 4577.050 3166.630 4579.120 ;
        RECT 0.000 4575.900 3165.930 4577.050 ;
        RECT 0.000 4574.645 3166.630 4575.900 ;
        RECT 0.000 4572.775 3165.930 4574.645 ;
        RECT 0.000 4571.710 3166.630 4572.775 ;
        RECT 0.700 4571.070 3166.630 4571.710 ;
        RECT 0.700 4570.560 3165.930 4571.070 ;
        RECT 0.000 4569.920 3165.930 4570.560 ;
        RECT 0.000 4568.490 3166.630 4569.920 ;
        RECT 0.700 4567.340 3166.630 4568.490 ;
        RECT 0.000 4565.270 3166.630 4567.340 ;
        RECT 0.700 4565.230 3166.630 4565.270 ;
        RECT 0.700 4564.120 3165.930 4565.230 ;
        RECT 0.000 4563.790 3165.930 4564.120 ;
        RECT 0.000 4562.510 3166.630 4563.790 ;
        RECT 0.700 4561.870 3166.630 4562.510 ;
        RECT 0.700 4561.360 3165.930 4561.870 ;
        RECT 0.000 4560.720 3165.930 4561.360 ;
        RECT 0.000 4552.670 3166.630 4560.720 ;
        RECT 0.000 4551.520 3165.930 4552.670 ;
        RECT 0.000 4533.920 3166.630 4551.520 ;
        RECT 0.700 4532.820 3166.630 4533.920 ;
        RECT 0.000 4523.920 3166.630 4532.820 ;
        RECT 0.700 4522.820 3166.630 4523.920 ;
        RECT 0.000 4424.420 3166.630 4522.820 ;
        RECT 0.700 4402.210 3166.630 4424.420 ;
        RECT 0.700 4401.810 3165.930 4402.210 ;
        RECT 0.700 4399.670 3122.620 4401.810 ;
        RECT 0.000 4398.980 3122.620 4399.670 ;
        RECT 0.700 4374.870 3122.620 4398.980 ;
        RECT 0.000 4374.220 3122.620 4374.870 ;
        RECT 0.700 4349.420 3122.620 4374.220 ;
        RECT 0.000 4327.610 3122.620 4349.420 ;
      LAYER met3 ;
        RECT 3122.620 4327.610 3167.855 4401.810 ;
      LAYER met3 ;
        RECT 0.000 4327.210 3165.930 4327.610 ;
        RECT 0.000 4213.010 3166.630 4327.210 ;
        RECT 0.700 4195.740 3166.630 4213.010 ;
        RECT 0.700 4194.630 3165.930 4195.740 ;
        RECT 0.700 4188.310 3166.630 4194.630 ;
        RECT 0.000 4185.740 3166.630 4188.310 ;
        RECT 0.000 4184.630 3165.930 4185.740 ;
        RECT 0.000 4180.270 3166.630 4184.630 ;
        RECT 0.000 4179.120 3165.930 4180.270 ;
        RECT 0.000 4177.510 3166.630 4179.120 ;
        RECT 0.000 4176.360 3165.930 4177.510 ;
        RECT 0.000 4174.290 3166.630 4176.360 ;
        RECT 0.000 4173.140 3165.930 4174.290 ;
        RECT 0.000 4171.070 3166.630 4173.140 ;
        RECT 0.000 4169.920 3165.930 4171.070 ;
        RECT 0.000 4163.110 3166.630 4169.920 ;
        RECT 0.700 4161.870 3166.630 4163.110 ;
        RECT 0.700 4160.720 3165.930 4161.870 ;
        RECT 0.700 4159.110 3166.630 4160.720 ;
        RECT 0.700 4157.960 3165.930 4159.110 ;
        RECT 0.700 4155.890 3166.630 4157.960 ;
        RECT 0.700 4154.740 3165.930 4155.890 ;
        RECT 0.700 4152.670 3166.630 4154.740 ;
        RECT 0.700 4151.520 3165.930 4152.670 ;
        RECT 0.700 4140.250 3166.630 4151.520 ;
        RECT 0.700 4139.100 3165.930 4140.250 ;
        RECT 0.700 4138.410 3166.630 4139.100 ;
        RECT 0.000 4137.490 3166.630 4138.410 ;
        RECT 0.000 4136.340 3165.930 4137.490 ;
        RECT 0.000 4134.270 3166.630 4136.340 ;
        RECT 0.000 4133.120 3165.930 4134.270 ;
        RECT 0.000 4131.050 3166.630 4133.120 ;
        RECT 0.000 4129.900 3165.930 4131.050 ;
        RECT 0.000 4128.645 3166.630 4129.900 ;
        RECT 0.000 4126.775 3165.930 4128.645 ;
        RECT 0.000 4125.070 3166.630 4126.775 ;
        RECT 0.000 4123.920 3165.930 4125.070 ;
        RECT 0.000 4119.230 3166.630 4123.920 ;
        RECT 0.000 4117.790 3165.930 4119.230 ;
        RECT 0.000 4115.870 3166.630 4117.790 ;
        RECT 0.000 4114.720 3165.930 4115.870 ;
        RECT 0.000 4106.670 3166.630 4114.720 ;
        RECT 0.000 4105.520 3165.930 4106.670 ;
        RECT 0.000 4002.010 3166.630 4105.520 ;
        RECT 0.700 3977.310 3166.630 4002.010 ;
        RECT 0.000 3956.220 3166.630 3977.310 ;
        RECT 0.000 3952.110 3165.930 3956.220 ;
        RECT 0.700 3931.520 3165.930 3952.110 ;
        RECT 0.700 3927.410 3166.630 3931.520 ;
        RECT 0.000 3906.330 3166.630 3927.410 ;
        RECT 0.000 3881.630 3165.930 3906.330 ;
        RECT 0.000 3787.110 3166.630 3881.630 ;
        RECT 0.700 3785.960 3166.630 3787.110 ;
        RECT 0.000 3777.910 3166.630 3785.960 ;
        RECT 0.700 3776.760 3166.630 3777.910 ;
        RECT 0.000 3774.840 3166.630 3776.760 ;
        RECT 0.700 3773.400 3166.630 3774.840 ;
        RECT 0.000 3768.710 3166.630 3773.400 ;
        RECT 0.700 3767.560 3166.630 3768.710 ;
        RECT 0.000 3765.855 3166.630 3767.560 ;
        RECT 0.700 3763.985 3166.630 3765.855 ;
        RECT 0.000 3762.730 3166.630 3763.985 ;
        RECT 0.700 3761.580 3166.630 3762.730 ;
        RECT 0.000 3759.510 3166.630 3761.580 ;
        RECT 0.700 3758.360 3166.630 3759.510 ;
        RECT 0.000 3756.290 3166.630 3758.360 ;
        RECT 0.700 3755.140 3166.630 3756.290 ;
        RECT 0.000 3753.530 3166.630 3755.140 ;
        RECT 0.700 3752.380 3166.630 3753.530 ;
        RECT 0.000 3750.740 3166.630 3752.380 ;
        RECT 0.000 3749.630 3165.930 3750.740 ;
        RECT 0.000 3741.110 3166.630 3749.630 ;
        RECT 0.700 3740.740 3166.630 3741.110 ;
        RECT 0.700 3739.960 3165.930 3740.740 ;
        RECT 0.000 3739.630 3165.930 3739.960 ;
        RECT 0.000 3737.890 3166.630 3739.630 ;
        RECT 0.700 3736.740 3166.630 3737.890 ;
        RECT 0.000 3734.670 3166.630 3736.740 ;
        RECT 0.700 3734.270 3166.630 3734.670 ;
        RECT 0.700 3733.520 3165.930 3734.270 ;
        RECT 0.000 3733.120 3165.930 3733.520 ;
        RECT 0.000 3731.910 3166.630 3733.120 ;
        RECT 0.700 3731.510 3166.630 3731.910 ;
        RECT 0.700 3730.760 3165.930 3731.510 ;
        RECT 0.000 3730.360 3165.930 3730.760 ;
        RECT 0.000 3728.290 3166.630 3730.360 ;
        RECT 0.000 3727.140 3165.930 3728.290 ;
        RECT 0.000 3725.070 3166.630 3727.140 ;
        RECT 0.000 3723.920 3165.930 3725.070 ;
        RECT 0.000 3722.710 3166.630 3723.920 ;
        RECT 0.700 3721.560 3166.630 3722.710 ;
        RECT 0.000 3719.490 3166.630 3721.560 ;
        RECT 0.700 3718.340 3166.630 3719.490 ;
        RECT 0.000 3716.270 3166.630 3718.340 ;
        RECT 0.700 3715.870 3166.630 3716.270 ;
        RECT 0.700 3715.120 3165.930 3715.870 ;
        RECT 0.000 3714.720 3165.930 3715.120 ;
        RECT 0.000 3713.510 3166.630 3714.720 ;
        RECT 0.700 3713.110 3166.630 3713.510 ;
        RECT 0.700 3712.360 3165.930 3713.110 ;
        RECT 0.000 3711.960 3165.930 3712.360 ;
        RECT 0.000 3709.890 3166.630 3711.960 ;
        RECT 0.000 3708.740 3165.930 3709.890 ;
        RECT 0.000 3706.670 3166.630 3708.740 ;
        RECT 0.000 3705.520 3165.930 3706.670 ;
        RECT 0.000 3694.250 3166.630 3705.520 ;
        RECT 0.000 3693.100 3165.930 3694.250 ;
        RECT 0.000 3691.490 3166.630 3693.100 ;
        RECT 0.000 3690.340 3165.930 3691.490 ;
        RECT 0.000 3688.270 3166.630 3690.340 ;
        RECT 0.000 3687.120 3165.930 3688.270 ;
        RECT 0.000 3685.050 3166.630 3687.120 ;
        RECT 0.000 3683.920 3165.930 3685.050 ;
        RECT 0.700 3683.900 3165.930 3683.920 ;
        RECT 0.700 3682.820 3166.630 3683.900 ;
        RECT 0.000 3682.645 3166.630 3682.820 ;
        RECT 0.000 3680.775 3165.930 3682.645 ;
        RECT 0.000 3679.070 3166.630 3680.775 ;
        RECT 0.000 3677.920 3165.930 3679.070 ;
        RECT 0.000 3673.920 3166.630 3677.920 ;
        RECT 0.700 3673.230 3166.630 3673.920 ;
        RECT 0.700 3672.820 3165.930 3673.230 ;
        RECT 0.000 3671.790 3165.930 3672.820 ;
        RECT 0.000 3669.870 3166.630 3671.790 ;
        RECT 0.000 3668.720 3165.930 3669.870 ;
        RECT 0.000 3660.670 3166.630 3668.720 ;
        RECT 0.000 3659.520 3165.930 3660.670 ;
        RECT 0.000 3571.110 3166.630 3659.520 ;
        RECT 0.700 3569.960 3166.630 3571.110 ;
        RECT 0.000 3561.910 3166.630 3569.960 ;
        RECT 0.700 3560.760 3166.630 3561.910 ;
        RECT 0.000 3558.840 3166.630 3560.760 ;
        RECT 0.700 3557.400 3166.630 3558.840 ;
        RECT 0.000 3552.710 3166.630 3557.400 ;
        RECT 0.700 3551.560 3166.630 3552.710 ;
        RECT 0.000 3549.855 3166.630 3551.560 ;
        RECT 0.700 3547.985 3166.630 3549.855 ;
        RECT 0.000 3546.730 3166.630 3547.985 ;
        RECT 0.700 3545.580 3166.630 3546.730 ;
        RECT 0.000 3543.510 3166.630 3545.580 ;
        RECT 0.700 3542.360 3166.630 3543.510 ;
        RECT 0.000 3540.290 3166.630 3542.360 ;
        RECT 0.700 3539.140 3166.630 3540.290 ;
        RECT 0.000 3537.530 3166.630 3539.140 ;
        RECT 0.700 3536.380 3166.630 3537.530 ;
        RECT 0.000 3525.740 3166.630 3536.380 ;
        RECT 0.000 3525.110 3165.930 3525.740 ;
        RECT 0.700 3524.630 3165.930 3525.110 ;
        RECT 0.700 3523.960 3166.630 3524.630 ;
        RECT 0.000 3521.890 3166.630 3523.960 ;
        RECT 0.700 3520.740 3166.630 3521.890 ;
        RECT 0.000 3518.670 3166.630 3520.740 ;
        RECT 0.700 3517.520 3166.630 3518.670 ;
        RECT 0.000 3515.910 3166.630 3517.520 ;
        RECT 0.700 3515.740 3166.630 3515.910 ;
        RECT 0.700 3514.760 3165.930 3515.740 ;
        RECT 0.000 3514.630 3165.930 3514.760 ;
        RECT 0.000 3509.270 3166.630 3514.630 ;
        RECT 0.000 3508.120 3165.930 3509.270 ;
        RECT 0.000 3506.710 3166.630 3508.120 ;
        RECT 0.700 3506.510 3166.630 3506.710 ;
        RECT 0.700 3505.560 3165.930 3506.510 ;
        RECT 0.000 3505.360 3165.930 3505.560 ;
        RECT 0.000 3503.490 3166.630 3505.360 ;
        RECT 0.700 3503.290 3166.630 3503.490 ;
        RECT 0.700 3502.340 3165.930 3503.290 ;
        RECT 0.000 3502.140 3165.930 3502.340 ;
        RECT 0.000 3500.270 3166.630 3502.140 ;
        RECT 0.700 3500.070 3166.630 3500.270 ;
        RECT 0.700 3499.120 3165.930 3500.070 ;
        RECT 0.000 3498.920 3165.930 3499.120 ;
        RECT 0.000 3497.510 3166.630 3498.920 ;
        RECT 0.700 3496.360 3166.630 3497.510 ;
        RECT 0.000 3490.870 3166.630 3496.360 ;
        RECT 0.000 3489.720 3165.930 3490.870 ;
        RECT 0.000 3488.110 3166.630 3489.720 ;
        RECT 0.000 3486.960 3165.930 3488.110 ;
        RECT 0.000 3484.890 3166.630 3486.960 ;
        RECT 0.000 3483.740 3165.930 3484.890 ;
        RECT 0.000 3481.670 3166.630 3483.740 ;
        RECT 0.000 3480.520 3165.930 3481.670 ;
        RECT 0.000 3469.250 3166.630 3480.520 ;
        RECT 0.000 3468.920 3165.930 3469.250 ;
        RECT 0.700 3468.100 3165.930 3468.920 ;
        RECT 0.700 3467.820 3166.630 3468.100 ;
        RECT 0.000 3466.490 3166.630 3467.820 ;
        RECT 0.000 3465.340 3165.930 3466.490 ;
        RECT 0.000 3463.270 3166.630 3465.340 ;
        RECT 0.000 3462.120 3165.930 3463.270 ;
        RECT 0.000 3460.050 3166.630 3462.120 ;
        RECT 0.000 3458.920 3165.930 3460.050 ;
        RECT 0.700 3458.900 3165.930 3458.920 ;
        RECT 0.700 3457.820 3166.630 3458.900 ;
        RECT 0.000 3457.645 3166.630 3457.820 ;
        RECT 0.000 3455.775 3165.930 3457.645 ;
        RECT 0.000 3454.070 3166.630 3455.775 ;
        RECT 0.000 3452.920 3165.930 3454.070 ;
        RECT 0.000 3448.230 3166.630 3452.920 ;
        RECT 0.000 3446.790 3165.930 3448.230 ;
        RECT 0.000 3444.870 3166.630 3446.790 ;
        RECT 0.000 3443.720 3165.930 3444.870 ;
        RECT 0.000 3435.670 3166.630 3443.720 ;
        RECT 0.000 3434.520 3165.930 3435.670 ;
        RECT 0.000 3355.110 3166.630 3434.520 ;
        RECT 0.700 3353.960 3166.630 3355.110 ;
        RECT 0.000 3345.910 3166.630 3353.960 ;
        RECT 0.700 3344.760 3166.630 3345.910 ;
        RECT 0.000 3342.840 3166.630 3344.760 ;
        RECT 0.700 3341.400 3166.630 3342.840 ;
        RECT 0.000 3336.710 3166.630 3341.400 ;
        RECT 0.700 3335.560 3166.630 3336.710 ;
        RECT 0.000 3333.855 3166.630 3335.560 ;
        RECT 0.700 3331.985 3166.630 3333.855 ;
        RECT 0.000 3330.730 3166.630 3331.985 ;
        RECT 0.700 3329.580 3166.630 3330.730 ;
        RECT 0.000 3327.510 3166.630 3329.580 ;
        RECT 0.700 3326.360 3166.630 3327.510 ;
        RECT 0.000 3324.290 3166.630 3326.360 ;
        RECT 0.700 3323.140 3166.630 3324.290 ;
        RECT 0.000 3321.530 3166.630 3323.140 ;
        RECT 0.700 3320.380 3166.630 3321.530 ;
        RECT 0.000 3309.110 3166.630 3320.380 ;
        RECT 0.700 3307.960 3166.630 3309.110 ;
        RECT 0.000 3305.890 3166.630 3307.960 ;
        RECT 0.700 3304.740 3166.630 3305.890 ;
        RECT 0.000 3302.670 3166.630 3304.740 ;
        RECT 0.700 3301.520 3166.630 3302.670 ;
        RECT 0.000 3300.740 3166.630 3301.520 ;
        RECT 0.000 3299.910 3165.930 3300.740 ;
        RECT 0.700 3299.630 3165.930 3299.910 ;
        RECT 0.700 3298.760 3166.630 3299.630 ;
        RECT 0.000 3290.740 3166.630 3298.760 ;
        RECT 0.000 3290.710 3165.930 3290.740 ;
        RECT 0.700 3289.630 3165.930 3290.710 ;
        RECT 0.700 3289.560 3166.630 3289.630 ;
        RECT 0.000 3287.490 3166.630 3289.560 ;
        RECT 0.700 3286.340 3166.630 3287.490 ;
        RECT 0.000 3284.270 3166.630 3286.340 ;
        RECT 0.700 3283.120 3165.930 3284.270 ;
        RECT 0.000 3281.510 3166.630 3283.120 ;
        RECT 0.700 3280.360 3165.930 3281.510 ;
        RECT 0.000 3278.290 3166.630 3280.360 ;
        RECT 0.000 3277.140 3165.930 3278.290 ;
        RECT 0.000 3275.070 3166.630 3277.140 ;
        RECT 0.000 3273.920 3165.930 3275.070 ;
        RECT 0.000 3265.870 3166.630 3273.920 ;
        RECT 0.000 3264.720 3165.930 3265.870 ;
        RECT 0.000 3263.110 3166.630 3264.720 ;
        RECT 0.000 3261.960 3165.930 3263.110 ;
        RECT 0.000 3259.890 3166.630 3261.960 ;
        RECT 0.000 3258.740 3165.930 3259.890 ;
        RECT 0.000 3256.670 3166.630 3258.740 ;
        RECT 0.000 3255.520 3165.930 3256.670 ;
        RECT 0.000 3253.920 3166.630 3255.520 ;
        RECT 0.700 3252.820 3166.630 3253.920 ;
        RECT 0.000 3244.250 3166.630 3252.820 ;
        RECT 0.000 3243.920 3165.930 3244.250 ;
        RECT 0.700 3243.100 3165.930 3243.920 ;
        RECT 0.700 3242.820 3166.630 3243.100 ;
        RECT 0.000 3241.490 3166.630 3242.820 ;
        RECT 0.000 3240.340 3165.930 3241.490 ;
        RECT 0.000 3238.270 3166.630 3240.340 ;
        RECT 0.000 3237.120 3165.930 3238.270 ;
        RECT 0.000 3235.050 3166.630 3237.120 ;
        RECT 0.000 3233.900 3165.930 3235.050 ;
        RECT 0.000 3232.645 3166.630 3233.900 ;
        RECT 0.000 3230.775 3165.930 3232.645 ;
        RECT 0.000 3229.070 3166.630 3230.775 ;
        RECT 0.000 3227.920 3165.930 3229.070 ;
        RECT 0.000 3223.230 3166.630 3227.920 ;
        RECT 0.000 3221.790 3165.930 3223.230 ;
        RECT 0.000 3219.870 3166.630 3221.790 ;
        RECT 0.000 3218.720 3165.930 3219.870 ;
        RECT 0.000 3210.670 3166.630 3218.720 ;
        RECT 0.000 3209.520 3165.930 3210.670 ;
        RECT 0.000 3139.110 3166.630 3209.520 ;
        RECT 0.700 3137.960 3166.630 3139.110 ;
        RECT 0.000 3129.910 3166.630 3137.960 ;
        RECT 0.700 3128.760 3166.630 3129.910 ;
        RECT 0.000 3126.840 3166.630 3128.760 ;
        RECT 0.700 3125.400 3166.630 3126.840 ;
        RECT 0.000 3120.710 3166.630 3125.400 ;
        RECT 0.700 3119.560 3166.630 3120.710 ;
        RECT 0.000 3117.855 3166.630 3119.560 ;
        RECT 0.700 3115.985 3166.630 3117.855 ;
        RECT 0.000 3114.730 3166.630 3115.985 ;
        RECT 0.700 3113.580 3166.630 3114.730 ;
        RECT 0.000 3111.510 3166.630 3113.580 ;
        RECT 0.700 3110.360 3166.630 3111.510 ;
        RECT 0.000 3108.290 3166.630 3110.360 ;
        RECT 0.700 3107.140 3166.630 3108.290 ;
        RECT 0.000 3105.530 3166.630 3107.140 ;
        RECT 0.700 3104.380 3166.630 3105.530 ;
        RECT 0.000 3093.110 3166.630 3104.380 ;
        RECT 0.700 3091.960 3166.630 3093.110 ;
        RECT 0.000 3089.890 3166.630 3091.960 ;
        RECT 0.700 3088.740 3166.630 3089.890 ;
        RECT 0.000 3086.670 3166.630 3088.740 ;
        RECT 0.700 3085.520 3166.630 3086.670 ;
        RECT 0.000 3083.910 3166.630 3085.520 ;
        RECT 0.700 3082.760 3166.630 3083.910 ;
        RECT 0.000 3075.740 3166.630 3082.760 ;
        RECT 0.000 3074.710 3165.930 3075.740 ;
        RECT 0.700 3074.630 3165.930 3074.710 ;
        RECT 0.700 3073.560 3166.630 3074.630 ;
        RECT 0.000 3071.490 3166.630 3073.560 ;
        RECT 0.700 3070.340 3166.630 3071.490 ;
        RECT 0.000 3068.270 3166.630 3070.340 ;
        RECT 0.700 3067.120 3166.630 3068.270 ;
        RECT 0.000 3065.740 3166.630 3067.120 ;
        RECT 0.000 3065.510 3165.930 3065.740 ;
        RECT 0.700 3064.630 3165.930 3065.510 ;
        RECT 0.700 3064.360 3166.630 3064.630 ;
        RECT 0.000 3058.270 3166.630 3064.360 ;
        RECT 0.000 3057.120 3165.930 3058.270 ;
        RECT 0.000 3055.510 3166.630 3057.120 ;
        RECT 0.000 3054.360 3165.930 3055.510 ;
        RECT 0.000 3052.290 3166.630 3054.360 ;
        RECT 0.000 3051.140 3165.930 3052.290 ;
        RECT 0.000 3049.070 3166.630 3051.140 ;
        RECT 0.000 3047.920 3165.930 3049.070 ;
        RECT 0.000 3039.870 3166.630 3047.920 ;
        RECT 0.000 3038.920 3165.930 3039.870 ;
        RECT 0.700 3038.720 3165.930 3038.920 ;
        RECT 0.700 3037.820 3166.630 3038.720 ;
        RECT 0.000 3037.110 3166.630 3037.820 ;
        RECT 0.000 3035.960 3165.930 3037.110 ;
        RECT 0.000 3033.890 3166.630 3035.960 ;
        RECT 0.000 3032.740 3165.930 3033.890 ;
        RECT 0.000 3030.670 3166.630 3032.740 ;
        RECT 0.000 3029.520 3165.930 3030.670 ;
        RECT 0.000 3028.920 3166.630 3029.520 ;
        RECT 0.700 3027.820 3166.630 3028.920 ;
        RECT 0.000 3018.250 3166.630 3027.820 ;
        RECT 0.000 3017.100 3165.930 3018.250 ;
        RECT 0.000 3015.490 3166.630 3017.100 ;
        RECT 0.000 3014.340 3165.930 3015.490 ;
        RECT 0.000 3012.270 3166.630 3014.340 ;
        RECT 0.000 3011.120 3165.930 3012.270 ;
        RECT 0.000 3009.050 3166.630 3011.120 ;
        RECT 0.000 3007.900 3165.930 3009.050 ;
        RECT 0.000 3006.645 3166.630 3007.900 ;
        RECT 0.000 3004.775 3165.930 3006.645 ;
        RECT 0.000 3003.070 3166.630 3004.775 ;
        RECT 0.000 3001.920 3165.930 3003.070 ;
        RECT 0.000 2997.230 3166.630 3001.920 ;
        RECT 0.000 2995.790 3165.930 2997.230 ;
        RECT 0.000 2993.870 3166.630 2995.790 ;
        RECT 0.000 2992.720 3165.930 2993.870 ;
        RECT 0.000 2984.670 3166.630 2992.720 ;
        RECT 0.000 2983.520 3165.930 2984.670 ;
        RECT 0.000 2923.110 3166.630 2983.520 ;
        RECT 0.700 2921.960 3166.630 2923.110 ;
        RECT 0.000 2913.910 3166.630 2921.960 ;
        RECT 0.700 2912.760 3166.630 2913.910 ;
        RECT 0.000 2910.840 3166.630 2912.760 ;
        RECT 0.700 2909.400 3166.630 2910.840 ;
        RECT 0.000 2904.710 3166.630 2909.400 ;
        RECT 0.700 2903.560 3166.630 2904.710 ;
        RECT 0.000 2901.855 3166.630 2903.560 ;
        RECT 0.700 2899.985 3166.630 2901.855 ;
        RECT 0.000 2898.730 3166.630 2899.985 ;
        RECT 0.700 2897.580 3166.630 2898.730 ;
        RECT 0.000 2895.510 3166.630 2897.580 ;
        RECT 0.700 2894.360 3166.630 2895.510 ;
        RECT 0.000 2892.290 3166.630 2894.360 ;
        RECT 0.700 2891.140 3166.630 2892.290 ;
        RECT 0.000 2889.530 3166.630 2891.140 ;
        RECT 0.700 2888.380 3166.630 2889.530 ;
        RECT 0.000 2877.110 3166.630 2888.380 ;
        RECT 0.700 2875.960 3166.630 2877.110 ;
        RECT 0.000 2873.890 3166.630 2875.960 ;
        RECT 0.700 2872.740 3166.630 2873.890 ;
        RECT 0.000 2870.670 3166.630 2872.740 ;
        RECT 0.700 2869.520 3166.630 2870.670 ;
        RECT 0.000 2867.910 3166.630 2869.520 ;
        RECT 0.700 2866.760 3166.630 2867.910 ;
        RECT 0.000 2858.710 3166.630 2866.760 ;
        RECT 0.700 2857.560 3166.630 2858.710 ;
        RECT 0.000 2855.490 3166.630 2857.560 ;
        RECT 0.700 2854.340 3166.630 2855.490 ;
        RECT 0.000 2852.270 3166.630 2854.340 ;
        RECT 0.700 2851.120 3166.630 2852.270 ;
        RECT 0.000 2850.740 3166.630 2851.120 ;
        RECT 0.000 2849.630 3165.930 2850.740 ;
        RECT 0.000 2849.510 3166.630 2849.630 ;
        RECT 0.700 2848.360 3166.630 2849.510 ;
        RECT 0.000 2840.740 3166.630 2848.360 ;
        RECT 0.000 2839.630 3165.930 2840.740 ;
        RECT 0.000 2833.270 3166.630 2839.630 ;
        RECT 0.000 2832.120 3165.930 2833.270 ;
        RECT 0.000 2830.510 3166.630 2832.120 ;
        RECT 0.000 2829.360 3165.930 2830.510 ;
        RECT 0.000 2827.290 3166.630 2829.360 ;
        RECT 0.000 2826.140 3165.930 2827.290 ;
        RECT 0.000 2824.070 3166.630 2826.140 ;
        RECT 0.000 2823.920 3165.930 2824.070 ;
        RECT 0.700 2822.920 3165.930 2823.920 ;
        RECT 0.700 2822.820 3166.630 2822.920 ;
        RECT 0.000 2814.870 3166.630 2822.820 ;
        RECT 0.000 2813.920 3165.930 2814.870 ;
        RECT 0.700 2813.720 3165.930 2813.920 ;
        RECT 0.700 2812.820 3166.630 2813.720 ;
        RECT 0.000 2812.110 3166.630 2812.820 ;
        RECT 0.000 2810.960 3165.930 2812.110 ;
        RECT 0.000 2808.890 3166.630 2810.960 ;
        RECT 0.000 2807.740 3165.930 2808.890 ;
        RECT 0.000 2805.670 3166.630 2807.740 ;
        RECT 0.000 2804.520 3165.930 2805.670 ;
        RECT 0.000 2793.250 3166.630 2804.520 ;
        RECT 0.000 2792.100 3165.930 2793.250 ;
        RECT 0.000 2790.490 3166.630 2792.100 ;
        RECT 0.000 2789.340 3165.930 2790.490 ;
        RECT 0.000 2787.270 3166.630 2789.340 ;
        RECT 0.000 2786.120 3165.930 2787.270 ;
        RECT 0.000 2784.050 3166.630 2786.120 ;
        RECT 0.000 2782.900 3165.930 2784.050 ;
        RECT 0.000 2781.645 3166.630 2782.900 ;
        RECT 0.000 2779.775 3165.930 2781.645 ;
        RECT 0.000 2778.070 3166.630 2779.775 ;
        RECT 0.000 2776.920 3165.930 2778.070 ;
        RECT 0.000 2772.230 3166.630 2776.920 ;
        RECT 0.000 2770.790 3165.930 2772.230 ;
        RECT 0.000 2768.870 3166.630 2770.790 ;
        RECT 0.000 2767.720 3165.930 2768.870 ;
        RECT 0.000 2759.670 3166.630 2767.720 ;
        RECT 0.000 2758.520 3165.930 2759.670 ;
        RECT 0.000 2707.110 3166.630 2758.520 ;
        RECT 0.700 2705.960 3166.630 2707.110 ;
        RECT 0.000 2697.910 3166.630 2705.960 ;
        RECT 0.700 2696.760 3166.630 2697.910 ;
        RECT 0.000 2694.840 3166.630 2696.760 ;
        RECT 0.700 2693.400 3166.630 2694.840 ;
        RECT 0.000 2688.710 3166.630 2693.400 ;
        RECT 0.700 2687.560 3166.630 2688.710 ;
        RECT 0.000 2685.855 3166.630 2687.560 ;
        RECT 0.700 2683.985 3166.630 2685.855 ;
        RECT 0.000 2682.730 3166.630 2683.985 ;
        RECT 0.700 2681.580 3166.630 2682.730 ;
        RECT 0.000 2679.510 3166.630 2681.580 ;
        RECT 0.700 2678.360 3166.630 2679.510 ;
        RECT 0.000 2676.290 3166.630 2678.360 ;
        RECT 0.700 2675.140 3166.630 2676.290 ;
        RECT 0.000 2673.530 3166.630 2675.140 ;
        RECT 0.700 2672.380 3166.630 2673.530 ;
        RECT 0.000 2661.110 3166.630 2672.380 ;
        RECT 0.700 2659.960 3166.630 2661.110 ;
        RECT 0.000 2657.890 3166.630 2659.960 ;
        RECT 0.700 2656.740 3166.630 2657.890 ;
        RECT 0.000 2654.670 3166.630 2656.740 ;
        RECT 0.700 2653.520 3166.630 2654.670 ;
        RECT 0.000 2651.910 3166.630 2653.520 ;
        RECT 0.700 2650.760 3166.630 2651.910 ;
        RECT 0.000 2642.710 3166.630 2650.760 ;
        RECT 0.700 2641.560 3166.630 2642.710 ;
        RECT 0.000 2639.490 3166.630 2641.560 ;
        RECT 0.700 2638.340 3166.630 2639.490 ;
        RECT 0.000 2636.270 3166.630 2638.340 ;
        RECT 0.700 2635.120 3166.630 2636.270 ;
        RECT 0.000 2633.510 3166.630 2635.120 ;
        RECT 0.700 2632.360 3166.630 2633.510 ;
        RECT 0.000 2625.740 3166.630 2632.360 ;
        RECT 0.000 2624.630 3165.930 2625.740 ;
        RECT 0.000 2615.735 3166.630 2624.630 ;
        RECT 0.000 2614.625 3165.930 2615.735 ;
        RECT 0.000 2608.920 3166.630 2614.625 ;
        RECT 0.700 2607.820 3166.630 2608.920 ;
        RECT 0.000 2607.270 3166.630 2607.820 ;
        RECT 0.000 2606.120 3165.930 2607.270 ;
        RECT 0.000 2604.510 3166.630 2606.120 ;
        RECT 0.000 2603.360 3165.930 2604.510 ;
        RECT 0.000 2601.290 3166.630 2603.360 ;
        RECT 0.000 2600.140 3165.930 2601.290 ;
        RECT 0.000 2598.920 3166.630 2600.140 ;
        RECT 0.700 2598.070 3166.630 2598.920 ;
        RECT 0.700 2597.820 3165.930 2598.070 ;
        RECT 0.000 2596.920 3165.930 2597.820 ;
        RECT 0.000 2588.870 3166.630 2596.920 ;
        RECT 0.000 2587.720 3165.930 2588.870 ;
        RECT 0.000 2586.110 3166.630 2587.720 ;
        RECT 0.000 2584.960 3165.930 2586.110 ;
        RECT 0.000 2582.890 3166.630 2584.960 ;
        RECT 0.000 2581.740 3165.930 2582.890 ;
        RECT 0.000 2579.670 3166.630 2581.740 ;
        RECT 0.000 2578.520 3165.930 2579.670 ;
        RECT 0.000 2567.250 3166.630 2578.520 ;
        RECT 0.000 2566.100 3165.930 2567.250 ;
        RECT 0.000 2564.490 3166.630 2566.100 ;
        RECT 0.000 2563.340 3165.930 2564.490 ;
        RECT 0.000 2561.270 3166.630 2563.340 ;
        RECT 0.000 2560.120 3165.930 2561.270 ;
        RECT 0.000 2558.050 3166.630 2560.120 ;
        RECT 0.000 2556.900 3165.930 2558.050 ;
        RECT 0.000 2555.645 3166.630 2556.900 ;
        RECT 0.000 2553.775 3165.930 2555.645 ;
        RECT 0.000 2552.070 3166.630 2553.775 ;
        RECT 0.000 2550.920 3165.930 2552.070 ;
        RECT 0.000 2546.230 3166.630 2550.920 ;
        RECT 0.000 2544.790 3165.930 2546.230 ;
        RECT 0.000 2542.870 3166.630 2544.790 ;
        RECT 0.000 2541.720 3165.930 2542.870 ;
        RECT 0.000 2533.670 3166.630 2541.720 ;
        RECT 0.000 2532.520 3165.930 2533.670 ;
        RECT 0.000 2491.110 3166.630 2532.520 ;
        RECT 0.700 2489.960 3166.630 2491.110 ;
        RECT 0.000 2481.910 3166.630 2489.960 ;
        RECT 0.700 2480.760 3166.630 2481.910 ;
        RECT 0.000 2478.840 3166.630 2480.760 ;
        RECT 0.700 2477.400 3166.630 2478.840 ;
        RECT 0.000 2472.710 3166.630 2477.400 ;
        RECT 0.700 2471.560 3166.630 2472.710 ;
        RECT 0.000 2469.855 3166.630 2471.560 ;
        RECT 0.700 2467.985 3166.630 2469.855 ;
        RECT 0.000 2466.730 3166.630 2467.985 ;
        RECT 0.700 2465.580 3166.630 2466.730 ;
        RECT 0.000 2463.510 3166.630 2465.580 ;
        RECT 0.700 2462.360 3166.630 2463.510 ;
        RECT 0.000 2460.290 3166.630 2462.360 ;
        RECT 0.700 2459.140 3166.630 2460.290 ;
        RECT 0.000 2457.530 3166.630 2459.140 ;
        RECT 0.700 2456.380 3166.630 2457.530 ;
        RECT 0.000 2445.110 3166.630 2456.380 ;
        RECT 0.700 2443.960 3166.630 2445.110 ;
        RECT 0.000 2441.890 3166.630 2443.960 ;
        RECT 0.700 2440.740 3166.630 2441.890 ;
        RECT 0.000 2438.670 3166.630 2440.740 ;
        RECT 0.700 2437.520 3166.630 2438.670 ;
        RECT 0.000 2435.910 3166.630 2437.520 ;
        RECT 0.700 2434.760 3166.630 2435.910 ;
        RECT 0.000 2426.710 3166.630 2434.760 ;
        RECT 0.700 2425.560 3166.630 2426.710 ;
        RECT 0.000 2423.490 3166.630 2425.560 ;
        RECT 0.700 2422.340 3166.630 2423.490 ;
        RECT 0.000 2420.270 3166.630 2422.340 ;
        RECT 0.700 2419.120 3166.630 2420.270 ;
        RECT 0.000 2417.510 3166.630 2419.120 ;
        RECT 0.700 2416.360 3166.630 2417.510 ;
        RECT 0.000 2393.920 3166.630 2416.360 ;
        RECT 0.700 2392.820 3166.630 2393.920 ;
        RECT 0.000 2383.920 3166.630 2392.820 ;
        RECT 0.700 2383.220 3166.630 2383.920 ;
        RECT 0.700 2382.820 3165.930 2383.220 ;
        RECT 0.000 2358.520 3165.930 2382.820 ;
        RECT 0.000 2333.320 3166.630 2358.520 ;
        RECT 0.000 2308.620 3165.930 2333.320 ;
        RECT 0.000 2279.000 3166.630 2308.620 ;
        RECT 0.700 2254.300 3166.630 2279.000 ;
        RECT 0.000 2229.110 3166.630 2254.300 ;
        RECT 0.700 2204.410 3166.630 2229.110 ;
        RECT 0.000 2163.210 3166.630 2204.410 ;
        RECT 0.000 2162.810 3165.930 2163.210 ;
        RECT 0.000 2088.610 3122.620 2162.810 ;
      LAYER met3 ;
        RECT 3122.620 2088.610 3167.855 2162.810 ;
      LAYER met3 ;
        RECT 0.000 2088.210 3165.930 2088.610 ;
        RECT 0.000 2068.420 3166.630 2088.210 ;
        RECT 0.700 2043.670 3166.630 2068.420 ;
        RECT 0.000 2042.970 3166.630 2043.670 ;
        RECT 0.700 2018.910 3166.630 2042.970 ;
        RECT 0.000 2018.210 3166.630 2018.910 ;
        RECT 0.700 1993.410 3166.630 2018.210 ;
        RECT 0.000 1942.220 3166.630 1993.410 ;
        RECT 0.000 1917.520 3165.930 1942.220 ;
        RECT 0.000 1892.330 3166.630 1917.520 ;
        RECT 0.000 1867.630 3165.930 1892.330 ;
        RECT 0.000 1853.110 3166.630 1867.630 ;
        RECT 0.700 1851.960 3166.630 1853.110 ;
        RECT 0.000 1843.910 3166.630 1851.960 ;
        RECT 0.700 1842.760 3166.630 1843.910 ;
        RECT 0.000 1840.840 3166.630 1842.760 ;
        RECT 0.700 1839.400 3166.630 1840.840 ;
        RECT 0.000 1834.710 3166.630 1839.400 ;
        RECT 0.700 1833.560 3166.630 1834.710 ;
        RECT 0.000 1831.855 3166.630 1833.560 ;
        RECT 0.700 1829.985 3166.630 1831.855 ;
        RECT 0.000 1828.730 3166.630 1829.985 ;
        RECT 0.700 1827.580 3166.630 1828.730 ;
        RECT 0.000 1825.510 3166.630 1827.580 ;
        RECT 0.700 1824.360 3166.630 1825.510 ;
        RECT 0.000 1822.290 3166.630 1824.360 ;
        RECT 0.700 1821.140 3166.630 1822.290 ;
        RECT 0.000 1819.530 3166.630 1821.140 ;
        RECT 0.700 1818.380 3166.630 1819.530 ;
        RECT 0.000 1807.110 3166.630 1818.380 ;
        RECT 0.700 1805.960 3166.630 1807.110 ;
        RECT 0.000 1803.890 3166.630 1805.960 ;
        RECT 0.700 1802.740 3166.630 1803.890 ;
        RECT 0.000 1800.670 3166.630 1802.740 ;
        RECT 0.700 1799.520 3166.630 1800.670 ;
        RECT 0.000 1797.910 3166.630 1799.520 ;
        RECT 0.700 1796.760 3166.630 1797.910 ;
        RECT 0.000 1788.710 3166.630 1796.760 ;
        RECT 0.700 1787.560 3166.630 1788.710 ;
        RECT 0.000 1785.490 3166.630 1787.560 ;
        RECT 0.700 1784.340 3166.630 1785.490 ;
        RECT 0.000 1782.270 3166.630 1784.340 ;
        RECT 0.700 1781.120 3166.630 1782.270 ;
        RECT 0.000 1779.510 3166.630 1781.120 ;
        RECT 0.700 1778.360 3166.630 1779.510 ;
        RECT 0.000 1748.920 3166.630 1778.360 ;
        RECT 0.700 1747.820 3166.630 1748.920 ;
        RECT 0.000 1740.740 3166.630 1747.820 ;
        RECT 0.000 1739.630 3165.930 1740.740 ;
        RECT 0.000 1738.920 3166.630 1739.630 ;
        RECT 0.700 1737.820 3166.630 1738.920 ;
        RECT 0.000 1730.735 3166.630 1737.820 ;
        RECT 0.000 1729.625 3165.930 1730.735 ;
        RECT 0.000 1721.270 3166.630 1729.625 ;
        RECT 0.000 1720.120 3165.930 1721.270 ;
        RECT 0.000 1718.510 3166.630 1720.120 ;
        RECT 0.000 1717.360 3165.930 1718.510 ;
        RECT 0.000 1715.290 3166.630 1717.360 ;
        RECT 0.000 1714.140 3165.930 1715.290 ;
        RECT 0.000 1712.070 3166.630 1714.140 ;
        RECT 0.000 1710.920 3165.930 1712.070 ;
        RECT 0.000 1702.870 3166.630 1710.920 ;
        RECT 0.000 1701.720 3165.930 1702.870 ;
        RECT 0.000 1700.110 3166.630 1701.720 ;
        RECT 0.000 1698.960 3165.930 1700.110 ;
        RECT 0.000 1696.890 3166.630 1698.960 ;
        RECT 0.000 1695.740 3165.930 1696.890 ;
        RECT 0.000 1693.670 3166.630 1695.740 ;
        RECT 0.000 1692.520 3165.930 1693.670 ;
        RECT 0.000 1681.250 3166.630 1692.520 ;
        RECT 0.000 1680.100 3165.930 1681.250 ;
        RECT 0.000 1678.490 3166.630 1680.100 ;
        RECT 0.000 1677.340 3165.930 1678.490 ;
        RECT 0.000 1675.270 3166.630 1677.340 ;
        RECT 0.000 1674.120 3165.930 1675.270 ;
        RECT 0.000 1672.050 3166.630 1674.120 ;
        RECT 0.000 1670.900 3165.930 1672.050 ;
        RECT 0.000 1669.645 3166.630 1670.900 ;
        RECT 0.000 1667.775 3165.930 1669.645 ;
        RECT 0.000 1666.070 3166.630 1667.775 ;
        RECT 0.000 1664.920 3165.930 1666.070 ;
        RECT 0.000 1660.230 3166.630 1664.920 ;
        RECT 0.000 1658.790 3165.930 1660.230 ;
        RECT 0.000 1656.870 3166.630 1658.790 ;
        RECT 0.000 1655.720 3165.930 1656.870 ;
        RECT 0.000 1647.670 3166.630 1655.720 ;
        RECT 0.000 1646.520 3165.930 1647.670 ;
        RECT 0.000 1637.110 3166.630 1646.520 ;
        RECT 0.700 1635.960 3166.630 1637.110 ;
        RECT 0.000 1627.910 3166.630 1635.960 ;
        RECT 0.700 1626.760 3166.630 1627.910 ;
        RECT 0.000 1624.840 3166.630 1626.760 ;
        RECT 0.700 1623.400 3166.630 1624.840 ;
        RECT 0.000 1618.710 3166.630 1623.400 ;
        RECT 0.700 1617.560 3166.630 1618.710 ;
        RECT 0.000 1615.855 3166.630 1617.560 ;
        RECT 0.700 1613.985 3166.630 1615.855 ;
        RECT 0.000 1612.730 3166.630 1613.985 ;
        RECT 0.700 1611.580 3166.630 1612.730 ;
        RECT 0.000 1609.510 3166.630 1611.580 ;
        RECT 0.700 1608.360 3166.630 1609.510 ;
        RECT 0.000 1606.290 3166.630 1608.360 ;
        RECT 0.700 1605.140 3166.630 1606.290 ;
        RECT 0.000 1603.530 3166.630 1605.140 ;
        RECT 0.700 1602.380 3166.630 1603.530 ;
        RECT 0.000 1591.110 3166.630 1602.380 ;
        RECT 0.700 1589.960 3166.630 1591.110 ;
        RECT 0.000 1587.890 3166.630 1589.960 ;
        RECT 0.700 1586.740 3166.630 1587.890 ;
        RECT 0.000 1584.670 3166.630 1586.740 ;
        RECT 0.700 1583.520 3166.630 1584.670 ;
        RECT 0.000 1581.910 3166.630 1583.520 ;
        RECT 0.700 1580.760 3166.630 1581.910 ;
        RECT 0.000 1572.710 3166.630 1580.760 ;
        RECT 0.700 1571.560 3166.630 1572.710 ;
        RECT 0.000 1569.490 3166.630 1571.560 ;
        RECT 0.700 1568.340 3166.630 1569.490 ;
        RECT 0.000 1566.270 3166.630 1568.340 ;
        RECT 0.700 1565.120 3166.630 1566.270 ;
        RECT 0.000 1563.510 3166.630 1565.120 ;
        RECT 0.700 1562.360 3166.630 1563.510 ;
        RECT 0.000 1533.920 3166.630 1562.360 ;
        RECT 0.700 1532.820 3166.630 1533.920 ;
        RECT 0.000 1523.920 3166.630 1532.820 ;
        RECT 0.700 1522.820 3166.630 1523.920 ;
        RECT 0.000 1515.740 3166.630 1522.820 ;
        RECT 0.000 1514.630 3165.930 1515.740 ;
        RECT 0.000 1505.735 3166.630 1514.630 ;
        RECT 0.000 1504.625 3165.930 1505.735 ;
        RECT 0.000 1495.270 3166.630 1504.625 ;
        RECT 0.000 1494.120 3165.930 1495.270 ;
        RECT 0.000 1492.510 3166.630 1494.120 ;
        RECT 0.000 1491.360 3165.930 1492.510 ;
        RECT 0.000 1489.290 3166.630 1491.360 ;
        RECT 0.000 1488.140 3165.930 1489.290 ;
        RECT 0.000 1486.070 3166.630 1488.140 ;
        RECT 0.000 1484.920 3165.930 1486.070 ;
        RECT 0.000 1476.870 3166.630 1484.920 ;
        RECT 0.000 1475.720 3165.930 1476.870 ;
        RECT 0.000 1474.110 3166.630 1475.720 ;
        RECT 0.000 1472.960 3165.930 1474.110 ;
        RECT 0.000 1470.890 3166.630 1472.960 ;
        RECT 0.000 1469.740 3165.930 1470.890 ;
        RECT 0.000 1467.670 3166.630 1469.740 ;
        RECT 0.000 1466.520 3165.930 1467.670 ;
        RECT 0.000 1455.250 3166.630 1466.520 ;
        RECT 0.000 1454.100 3165.930 1455.250 ;
        RECT 0.000 1452.490 3166.630 1454.100 ;
        RECT 0.000 1451.340 3165.930 1452.490 ;
        RECT 0.000 1449.270 3166.630 1451.340 ;
        RECT 0.000 1448.120 3165.930 1449.270 ;
        RECT 0.000 1446.050 3166.630 1448.120 ;
        RECT 0.000 1444.900 3165.930 1446.050 ;
        RECT 0.000 1443.645 3166.630 1444.900 ;
        RECT 0.000 1441.775 3165.930 1443.645 ;
        RECT 0.000 1440.070 3166.630 1441.775 ;
        RECT 0.000 1438.920 3165.930 1440.070 ;
        RECT 0.000 1434.230 3166.630 1438.920 ;
        RECT 0.000 1432.790 3165.930 1434.230 ;
        RECT 0.000 1430.870 3166.630 1432.790 ;
        RECT 0.000 1429.720 3165.930 1430.870 ;
        RECT 0.000 1421.670 3166.630 1429.720 ;
        RECT 0.000 1421.110 3165.930 1421.670 ;
        RECT 0.700 1420.520 3165.930 1421.110 ;
        RECT 0.700 1419.960 3166.630 1420.520 ;
        RECT 0.000 1411.910 3166.630 1419.960 ;
        RECT 0.700 1410.760 3166.630 1411.910 ;
        RECT 0.000 1408.840 3166.630 1410.760 ;
        RECT 0.700 1407.400 3166.630 1408.840 ;
        RECT 0.000 1402.710 3166.630 1407.400 ;
        RECT 0.700 1401.560 3166.630 1402.710 ;
        RECT 0.000 1399.855 3166.630 1401.560 ;
        RECT 0.700 1397.985 3166.630 1399.855 ;
        RECT 0.000 1396.730 3166.630 1397.985 ;
        RECT 0.700 1395.580 3166.630 1396.730 ;
        RECT 0.000 1393.510 3166.630 1395.580 ;
        RECT 0.700 1392.360 3166.630 1393.510 ;
        RECT 0.000 1390.290 3166.630 1392.360 ;
        RECT 0.700 1389.140 3166.630 1390.290 ;
        RECT 0.000 1387.530 3166.630 1389.140 ;
        RECT 0.700 1386.380 3166.630 1387.530 ;
        RECT 0.000 1375.110 3166.630 1386.380 ;
        RECT 0.700 1373.960 3166.630 1375.110 ;
        RECT 0.000 1371.890 3166.630 1373.960 ;
        RECT 0.700 1370.740 3166.630 1371.890 ;
        RECT 0.000 1368.670 3166.630 1370.740 ;
        RECT 0.700 1367.520 3166.630 1368.670 ;
        RECT 0.000 1365.910 3166.630 1367.520 ;
        RECT 0.700 1364.760 3166.630 1365.910 ;
        RECT 0.000 1356.710 3166.630 1364.760 ;
        RECT 0.700 1355.560 3166.630 1356.710 ;
        RECT 0.000 1353.490 3166.630 1355.560 ;
        RECT 0.700 1352.340 3166.630 1353.490 ;
        RECT 0.000 1350.270 3166.630 1352.340 ;
        RECT 0.700 1349.120 3166.630 1350.270 ;
        RECT 0.000 1347.510 3166.630 1349.120 ;
        RECT 0.700 1346.360 3166.630 1347.510 ;
        RECT 0.000 1318.920 3166.630 1346.360 ;
        RECT 0.700 1317.820 3166.630 1318.920 ;
        RECT 0.000 1308.920 3166.630 1317.820 ;
        RECT 0.700 1307.820 3166.630 1308.920 ;
        RECT 0.000 1290.740 3166.630 1307.820 ;
        RECT 0.000 1289.630 3165.930 1290.740 ;
        RECT 0.000 1280.735 3166.630 1289.630 ;
        RECT 0.000 1279.625 3165.930 1280.735 ;
        RECT 0.000 1270.270 3166.630 1279.625 ;
        RECT 0.000 1269.120 3165.930 1270.270 ;
        RECT 0.000 1267.510 3166.630 1269.120 ;
        RECT 0.000 1266.360 3165.930 1267.510 ;
        RECT 0.000 1264.290 3166.630 1266.360 ;
        RECT 0.000 1263.140 3165.930 1264.290 ;
        RECT 0.000 1261.070 3166.630 1263.140 ;
        RECT 0.000 1259.920 3165.930 1261.070 ;
        RECT 0.000 1251.870 3166.630 1259.920 ;
        RECT 0.000 1250.720 3165.930 1251.870 ;
        RECT 0.000 1249.110 3166.630 1250.720 ;
        RECT 0.000 1247.960 3165.930 1249.110 ;
        RECT 0.000 1245.890 3166.630 1247.960 ;
        RECT 0.000 1244.740 3165.930 1245.890 ;
        RECT 0.000 1242.670 3166.630 1244.740 ;
        RECT 0.000 1241.520 3165.930 1242.670 ;
        RECT 0.000 1230.250 3166.630 1241.520 ;
        RECT 0.000 1229.100 3165.930 1230.250 ;
        RECT 0.000 1227.490 3166.630 1229.100 ;
        RECT 0.000 1226.340 3165.930 1227.490 ;
        RECT 0.000 1224.270 3166.630 1226.340 ;
        RECT 0.000 1223.120 3165.930 1224.270 ;
        RECT 0.000 1221.050 3166.630 1223.120 ;
        RECT 0.000 1219.900 3165.930 1221.050 ;
        RECT 0.000 1218.645 3166.630 1219.900 ;
        RECT 0.000 1216.775 3165.930 1218.645 ;
        RECT 0.000 1215.070 3166.630 1216.775 ;
        RECT 0.000 1213.920 3165.930 1215.070 ;
        RECT 0.000 1209.230 3166.630 1213.920 ;
        RECT 0.000 1207.790 3165.930 1209.230 ;
        RECT 0.000 1205.870 3166.630 1207.790 ;
        RECT 0.000 1205.110 3165.930 1205.870 ;
        RECT 0.700 1204.720 3165.930 1205.110 ;
        RECT 0.700 1203.960 3166.630 1204.720 ;
        RECT 0.000 1196.670 3166.630 1203.960 ;
        RECT 0.000 1195.910 3165.930 1196.670 ;
        RECT 0.700 1195.520 3165.930 1195.910 ;
        RECT 0.700 1194.760 3166.630 1195.520 ;
        RECT 0.000 1192.840 3166.630 1194.760 ;
        RECT 0.700 1191.400 3166.630 1192.840 ;
        RECT 0.000 1186.710 3166.630 1191.400 ;
        RECT 0.700 1185.560 3166.630 1186.710 ;
        RECT 0.000 1183.855 3166.630 1185.560 ;
        RECT 0.700 1181.985 3166.630 1183.855 ;
        RECT 0.000 1180.730 3166.630 1181.985 ;
        RECT 0.700 1179.580 3166.630 1180.730 ;
        RECT 0.000 1177.510 3166.630 1179.580 ;
        RECT 0.700 1176.360 3166.630 1177.510 ;
        RECT 0.000 1174.290 3166.630 1176.360 ;
        RECT 0.700 1173.140 3166.630 1174.290 ;
        RECT 0.000 1171.530 3166.630 1173.140 ;
        RECT 0.700 1170.380 3166.630 1171.530 ;
        RECT 0.000 1159.110 3166.630 1170.380 ;
        RECT 0.700 1157.960 3166.630 1159.110 ;
        RECT 0.000 1155.890 3166.630 1157.960 ;
        RECT 0.700 1154.740 3166.630 1155.890 ;
        RECT 0.000 1152.670 3166.630 1154.740 ;
        RECT 0.700 1151.520 3166.630 1152.670 ;
        RECT 0.000 1149.910 3166.630 1151.520 ;
        RECT 0.700 1148.760 3166.630 1149.910 ;
        RECT 0.000 1140.710 3166.630 1148.760 ;
        RECT 0.700 1139.560 3166.630 1140.710 ;
        RECT 0.000 1137.490 3166.630 1139.560 ;
        RECT 0.700 1136.340 3166.630 1137.490 ;
        RECT 0.000 1134.270 3166.630 1136.340 ;
        RECT 0.700 1133.120 3166.630 1134.270 ;
        RECT 0.000 1131.510 3166.630 1133.120 ;
        RECT 0.700 1130.360 3166.630 1131.510 ;
        RECT 0.000 1103.920 3166.630 1130.360 ;
        RECT 0.700 1102.820 3166.630 1103.920 ;
        RECT 0.000 1093.920 3166.630 1102.820 ;
        RECT 0.700 1092.820 3166.630 1093.920 ;
        RECT 0.000 1065.740 3166.630 1092.820 ;
        RECT 0.000 1064.630 3165.930 1065.740 ;
        RECT 0.000 1055.735 3166.630 1064.630 ;
        RECT 0.000 1054.625 3165.930 1055.735 ;
        RECT 0.000 1045.270 3166.630 1054.625 ;
        RECT 0.000 1044.120 3165.930 1045.270 ;
        RECT 0.000 1042.510 3166.630 1044.120 ;
        RECT 0.000 1041.360 3165.930 1042.510 ;
        RECT 0.000 1039.290 3166.630 1041.360 ;
        RECT 0.000 1038.140 3165.930 1039.290 ;
        RECT 0.000 1036.070 3166.630 1038.140 ;
        RECT 0.000 1034.920 3165.930 1036.070 ;
        RECT 0.000 1026.870 3166.630 1034.920 ;
        RECT 0.000 1025.720 3165.930 1026.870 ;
        RECT 0.000 1024.110 3166.630 1025.720 ;
        RECT 0.000 1022.960 3165.930 1024.110 ;
        RECT 0.000 1020.890 3166.630 1022.960 ;
        RECT 0.000 1019.740 3165.930 1020.890 ;
        RECT 0.000 1017.670 3166.630 1019.740 ;
        RECT 0.000 1016.520 3165.930 1017.670 ;
        RECT 0.000 1005.250 3166.630 1016.520 ;
        RECT 0.000 1004.100 3165.930 1005.250 ;
        RECT 0.000 1002.490 3166.630 1004.100 ;
        RECT 0.000 1001.340 3165.930 1002.490 ;
        RECT 0.000 999.270 3166.630 1001.340 ;
        RECT 0.000 998.120 3165.930 999.270 ;
        RECT 0.000 996.050 3166.630 998.120 ;
        RECT 0.000 994.900 3165.930 996.050 ;
        RECT 0.000 993.645 3166.630 994.900 ;
        RECT 0.000 991.775 3165.930 993.645 ;
        RECT 0.000 990.070 3166.630 991.775 ;
        RECT 0.000 989.110 3165.930 990.070 ;
        RECT 0.700 988.920 3165.930 989.110 ;
        RECT 0.700 987.960 3166.630 988.920 ;
        RECT 0.000 984.230 3166.630 987.960 ;
        RECT 0.000 982.790 3165.930 984.230 ;
        RECT 0.000 980.870 3166.630 982.790 ;
        RECT 0.000 979.910 3165.930 980.870 ;
        RECT 0.700 979.720 3165.930 979.910 ;
        RECT 0.700 978.760 3166.630 979.720 ;
        RECT 0.000 976.840 3166.630 978.760 ;
        RECT 0.700 975.400 3166.630 976.840 ;
        RECT 0.000 971.670 3166.630 975.400 ;
        RECT 0.000 970.710 3165.930 971.670 ;
        RECT 0.700 970.520 3165.930 970.710 ;
        RECT 0.700 969.560 3166.630 970.520 ;
        RECT 0.000 967.855 3166.630 969.560 ;
        RECT 0.700 965.985 3166.630 967.855 ;
        RECT 0.000 964.730 3166.630 965.985 ;
        RECT 0.700 963.580 3166.630 964.730 ;
        RECT 0.000 961.510 3166.630 963.580 ;
        RECT 0.700 960.360 3166.630 961.510 ;
        RECT 0.000 958.290 3166.630 960.360 ;
        RECT 0.700 957.140 3166.630 958.290 ;
        RECT 0.000 955.530 3166.630 957.140 ;
        RECT 0.700 954.380 3166.630 955.530 ;
        RECT 0.000 943.110 3166.630 954.380 ;
        RECT 0.700 941.960 3166.630 943.110 ;
        RECT 0.000 939.890 3166.630 941.960 ;
        RECT 0.700 938.740 3166.630 939.890 ;
        RECT 0.000 936.670 3166.630 938.740 ;
        RECT 0.700 935.520 3166.630 936.670 ;
        RECT 0.000 933.910 3166.630 935.520 ;
        RECT 0.700 932.760 3166.630 933.910 ;
        RECT 0.000 924.710 3166.630 932.760 ;
        RECT 0.700 923.560 3166.630 924.710 ;
        RECT 0.000 921.490 3166.630 923.560 ;
        RECT 0.700 920.340 3166.630 921.490 ;
        RECT 0.000 918.270 3166.630 920.340 ;
        RECT 0.700 917.120 3166.630 918.270 ;
        RECT 0.000 915.510 3166.630 917.120 ;
        RECT 0.700 914.360 3166.630 915.510 ;
        RECT 0.000 888.920 3166.630 914.360 ;
        RECT 0.700 887.820 3166.630 888.920 ;
        RECT 0.000 878.920 3166.630 887.820 ;
        RECT 0.700 877.820 3166.630 878.920 ;
        RECT 0.000 840.740 3166.630 877.820 ;
        RECT 0.000 839.630 3165.930 840.740 ;
        RECT 0.000 830.735 3166.630 839.630 ;
        RECT 0.000 829.625 3165.930 830.735 ;
        RECT 0.000 819.270 3166.630 829.625 ;
        RECT 0.000 818.120 3165.930 819.270 ;
        RECT 0.000 816.510 3166.630 818.120 ;
        RECT 0.000 815.360 3165.930 816.510 ;
        RECT 0.000 813.290 3166.630 815.360 ;
        RECT 0.000 812.140 3165.930 813.290 ;
        RECT 0.000 810.070 3166.630 812.140 ;
        RECT 0.000 808.920 3165.930 810.070 ;
        RECT 0.000 800.870 3166.630 808.920 ;
        RECT 0.000 799.720 3165.930 800.870 ;
        RECT 0.000 798.110 3166.630 799.720 ;
        RECT 0.000 796.960 3165.930 798.110 ;
        RECT 0.000 794.890 3166.630 796.960 ;
        RECT 0.000 793.740 3165.930 794.890 ;
        RECT 0.000 791.670 3166.630 793.740 ;
        RECT 0.000 790.520 3165.930 791.670 ;
        RECT 0.000 779.250 3166.630 790.520 ;
        RECT 0.000 778.100 3165.930 779.250 ;
        RECT 0.000 776.490 3166.630 778.100 ;
        RECT 0.000 775.340 3165.930 776.490 ;
        RECT 0.000 773.270 3166.630 775.340 ;
        RECT 0.000 773.110 3165.930 773.270 ;
        RECT 0.700 772.120 3165.930 773.110 ;
        RECT 0.700 771.960 3166.630 772.120 ;
        RECT 0.000 770.050 3166.630 771.960 ;
        RECT 0.000 768.900 3165.930 770.050 ;
        RECT 0.000 767.645 3166.630 768.900 ;
        RECT 0.000 765.775 3165.930 767.645 ;
        RECT 0.000 764.070 3166.630 765.775 ;
        RECT 0.000 763.910 3165.930 764.070 ;
        RECT 0.700 762.920 3165.930 763.910 ;
        RECT 0.700 762.760 3166.630 762.920 ;
        RECT 0.000 760.840 3166.630 762.760 ;
        RECT 0.700 759.400 3166.630 760.840 ;
        RECT 0.000 758.230 3166.630 759.400 ;
        RECT 0.000 756.790 3165.930 758.230 ;
        RECT 0.000 754.870 3166.630 756.790 ;
        RECT 0.000 754.710 3165.930 754.870 ;
        RECT 0.700 753.720 3165.930 754.710 ;
        RECT 0.700 753.560 3166.630 753.720 ;
        RECT 0.000 751.855 3166.630 753.560 ;
        RECT 0.700 749.985 3166.630 751.855 ;
        RECT 0.000 748.730 3166.630 749.985 ;
        RECT 0.700 747.580 3166.630 748.730 ;
        RECT 0.000 745.670 3166.630 747.580 ;
        RECT 0.000 745.510 3165.930 745.670 ;
        RECT 0.700 744.520 3165.930 745.510 ;
        RECT 0.700 744.360 3166.630 744.520 ;
        RECT 0.000 742.290 3166.630 744.360 ;
        RECT 0.700 741.140 3166.630 742.290 ;
        RECT 0.000 739.530 3166.630 741.140 ;
        RECT 0.700 738.380 3166.630 739.530 ;
        RECT 0.000 727.110 3166.630 738.380 ;
        RECT 0.700 725.960 3166.630 727.110 ;
        RECT 0.000 723.890 3166.630 725.960 ;
        RECT 0.700 722.740 3166.630 723.890 ;
        RECT 0.000 720.670 3166.630 722.740 ;
        RECT 0.700 719.520 3166.630 720.670 ;
        RECT 0.000 717.910 3166.630 719.520 ;
        RECT 0.700 716.760 3166.630 717.910 ;
        RECT 0.000 708.710 3166.630 716.760 ;
        RECT 0.700 707.560 3166.630 708.710 ;
        RECT 0.000 705.490 3166.630 707.560 ;
        RECT 0.700 704.340 3166.630 705.490 ;
        RECT 0.000 702.270 3166.630 704.340 ;
        RECT 0.700 701.120 3166.630 702.270 ;
        RECT 0.000 699.510 3166.630 701.120 ;
        RECT 0.700 698.360 3166.630 699.510 ;
        RECT 0.000 673.920 3166.630 698.360 ;
        RECT 0.700 672.820 3166.630 673.920 ;
        RECT 0.000 663.920 3166.630 672.820 ;
        RECT 0.700 662.820 3166.630 663.920 ;
        RECT 0.000 615.740 3166.630 662.820 ;
        RECT 0.000 614.630 3165.930 615.740 ;
        RECT 0.000 605.735 3166.630 614.630 ;
        RECT 0.000 604.625 3165.930 605.735 ;
        RECT 0.000 594.270 3166.630 604.625 ;
        RECT 0.000 593.120 3165.930 594.270 ;
        RECT 0.000 591.510 3166.630 593.120 ;
        RECT 0.000 590.360 3165.930 591.510 ;
        RECT 0.000 588.290 3166.630 590.360 ;
        RECT 0.000 587.140 3165.930 588.290 ;
        RECT 0.000 585.070 3166.630 587.140 ;
        RECT 0.000 583.920 3165.930 585.070 ;
        RECT 0.000 575.870 3166.630 583.920 ;
        RECT 0.000 574.720 3165.930 575.870 ;
        RECT 0.000 573.110 3166.630 574.720 ;
        RECT 0.000 571.960 3165.930 573.110 ;
        RECT 0.000 569.890 3166.630 571.960 ;
        RECT 0.000 568.740 3165.930 569.890 ;
        RECT 0.000 566.670 3166.630 568.740 ;
        RECT 0.000 565.520 3165.930 566.670 ;
        RECT 0.000 554.250 3166.630 565.520 ;
        RECT 0.000 553.100 3165.930 554.250 ;
        RECT 0.000 551.490 3166.630 553.100 ;
        RECT 0.000 550.340 3165.930 551.490 ;
        RECT 0.000 548.270 3166.630 550.340 ;
        RECT 0.000 547.120 3165.930 548.270 ;
        RECT 0.000 545.050 3166.630 547.120 ;
        RECT 0.000 543.900 3165.930 545.050 ;
        RECT 0.000 542.645 3166.630 543.900 ;
        RECT 0.000 540.775 3165.930 542.645 ;
        RECT 0.000 539.070 3166.630 540.775 ;
        RECT 0.000 537.920 3165.930 539.070 ;
        RECT 0.000 533.230 3166.630 537.920 ;
        RECT 0.000 531.790 3165.930 533.230 ;
        RECT 0.000 529.870 3166.630 531.790 ;
        RECT 0.000 528.720 3165.930 529.870 ;
        RECT 0.000 520.670 3166.630 528.720 ;
        RECT 0.000 519.520 3165.930 520.670 ;
        RECT 0.000 415.000 3166.630 519.520 ;
        RECT 0.700 390.740 3166.630 415.000 ;
        RECT 0.700 390.300 3165.930 390.740 ;
        RECT 0.000 389.630 3165.930 390.300 ;
        RECT 0.000 380.735 3166.630 389.630 ;
        RECT 0.000 379.625 3165.930 380.735 ;
        RECT 0.000 368.270 3166.630 379.625 ;
        RECT 0.000 367.120 3165.930 368.270 ;
        RECT 0.000 365.510 3166.630 367.120 ;
        RECT 0.000 365.110 3165.930 365.510 ;
        RECT 0.700 364.360 3165.930 365.110 ;
        RECT 0.700 362.290 3166.630 364.360 ;
        RECT 0.700 361.140 3165.930 362.290 ;
        RECT 0.700 359.070 3166.630 361.140 ;
        RECT 0.700 357.920 3165.930 359.070 ;
        RECT 0.700 349.870 3166.630 357.920 ;
        RECT 0.700 348.720 3165.930 349.870 ;
        RECT 0.700 347.110 3166.630 348.720 ;
        RECT 0.700 345.960 3165.930 347.110 ;
        RECT 0.700 343.890 3166.630 345.960 ;
        RECT 0.700 342.740 3165.930 343.890 ;
        RECT 0.700 340.670 3166.630 342.740 ;
        RECT 0.700 340.410 3165.930 340.670 ;
        RECT 0.000 339.520 3165.930 340.410 ;
        RECT 0.000 328.250 3166.630 339.520 ;
        RECT 0.000 327.100 3165.930 328.250 ;
        RECT 0.000 325.490 3166.630 327.100 ;
        RECT 0.000 324.340 3165.930 325.490 ;
        RECT 0.000 322.270 3166.630 324.340 ;
        RECT 0.000 321.120 3165.930 322.270 ;
        RECT 0.000 319.050 3166.630 321.120 ;
        RECT 0.000 317.900 3165.930 319.050 ;
        RECT 0.000 316.645 3166.630 317.900 ;
        RECT 0.000 314.775 3165.930 316.645 ;
        RECT 0.000 313.070 3166.630 314.775 ;
        RECT 0.000 311.920 3165.930 313.070 ;
        RECT 0.000 307.230 3166.630 311.920 ;
        RECT 0.000 305.790 3165.930 307.230 ;
        RECT 0.000 303.870 3166.630 305.790 ;
        RECT 0.000 302.720 3165.930 303.870 ;
        RECT 0.000 294.670 3166.630 302.720 ;
        RECT 0.000 293.520 3165.930 294.670 ;
        RECT 0.000 268.725 3166.630 293.520 ;
        RECT 0.700 265.335 3166.630 268.725 ;
        RECT 0.000 204.420 3166.630 265.335 ;
        RECT 0.700 179.670 3166.630 204.420 ;
        RECT 0.000 154.210 3166.630 179.670 ;
        RECT 0.700 129.410 3166.630 154.210 ;
        RECT 0.000 13.775 3166.630 129.410 ;
      LAYER met4 ;
        RECT 2873.760 245.640 2894.850 3722.280 ;
        RECT 2902.050 245.640 2904.450 3722.280 ;
        RECT 2911.650 245.640 2934.850 3722.280 ;
        RECT 2942.050 245.640 2974.850 3722.280 ;
        RECT 2982.050 245.640 2984.450 3722.280 ;
        RECT 2991.650 2213.045 3014.850 3722.280 ;
        RECT 3022.050 2213.045 3034.065 3722.280 ;
        RECT 2991.650 1472.675 3034.065 2213.045 ;
        RECT 2991.650 245.640 3014.850 1472.675 ;
        RECT 3022.050 245.640 3034.065 1472.675 ;
  END
END openframe_project_wrapper
END LIBRARY

